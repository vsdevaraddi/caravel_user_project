magic
tech sky130A
magscale 1 2
timestamp 1647698485
<< checkpaint >>
rect -12658 -11586 596582 715522
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 328454 700952 328460 701004
rect 328512 700992 328518 701004
rect 413646 700992 413652 701004
rect 328512 700964 413652 700992
rect 328512 700952 328518 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 218974 700884 218980 700936
rect 219032 700924 219038 700936
rect 338758 700924 338764 700936
rect 219032 700896 338764 700924
rect 219032 700884 219038 700896
rect 338758 700884 338764 700896
rect 338816 700884 338822 700936
rect 202782 700816 202788 700868
rect 202840 700856 202846 700868
rect 337378 700856 337384 700868
rect 202840 700828 337384 700856
rect 202840 700816 202846 700828
rect 337378 700816 337384 700828
rect 337436 700816 337442 700868
rect 322934 700748 322940 700800
rect 322992 700788 322998 700800
rect 478506 700788 478512 700800
rect 322992 700760 478512 700788
rect 322992 700748 322998 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 154114 700680 154120 700732
rect 154172 700720 154178 700732
rect 344278 700720 344284 700732
rect 154172 700692 344284 700720
rect 154172 700680 154178 700692
rect 344278 700680 344284 700692
rect 344336 700680 344342 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 342898 700652 342904 700664
rect 137888 700624 342904 700652
rect 137888 700612 137894 700624
rect 342898 700612 342904 700624
rect 342956 700612 342962 700664
rect 317414 700544 317420 700596
rect 317472 700584 317478 700596
rect 543458 700584 543464 700596
rect 317472 700556 543464 700584
rect 317472 700544 317478 700556
rect 543458 700544 543464 700556
rect 543516 700544 543522 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 349798 700516 349804 700528
rect 89220 700488 349804 700516
rect 89220 700476 89226 700488
rect 349798 700476 349804 700488
rect 349856 700476 349862 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 348418 700448 348424 700460
rect 73028 700420 348424 700448
rect 73028 700408 73034 700420
rect 348418 700408 348424 700420
rect 348476 700408 348482 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 355318 700380 355324 700392
rect 24360 700352 355324 700380
rect 24360 700340 24366 700352
rect 355318 700340 355324 700352
rect 355376 700340 355382 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 353938 700312 353944 700324
rect 8168 700284 353944 700312
rect 8168 700272 8174 700284
rect 353938 700272 353944 700284
rect 353996 700272 354002 700324
rect 325694 700204 325700 700256
rect 325752 700244 325758 700256
rect 397454 700244 397460 700256
rect 325752 700216 397460 700244
rect 325752 700204 325758 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 267642 700136 267648 700188
rect 267700 700176 267706 700188
rect 335998 700176 336004 700188
rect 267700 700148 336004 700176
rect 267700 700136 267706 700148
rect 335998 700136 336004 700148
rect 336056 700136 336062 700188
rect 333974 700068 333980 700120
rect 334032 700108 334038 700120
rect 348786 700108 348792 700120
rect 334032 700080 348792 700108
rect 334032 700068 334038 700080
rect 348786 700068 348792 700080
rect 348844 700068 348850 700120
rect 310514 696940 310520 696992
rect 310572 696980 310578 696992
rect 580166 696980 580172 696992
rect 310572 696952 580172 696980
rect 310572 696940 310578 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 311894 683204 311900 683256
rect 311952 683244 311958 683256
rect 580166 683244 580172 683256
rect 311952 683216 580172 683244
rect 311952 683204 311958 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 361574 683176 361580 683188
rect 3476 683148 361580 683176
rect 3476 683136 3482 683148
rect 361574 683136 361580 683148
rect 361632 683136 361638 683188
rect 309134 670760 309140 670812
rect 309192 670800 309198 670812
rect 580166 670800 580172 670812
rect 309192 670772 580172 670800
rect 309192 670760 309198 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 364426 670732 364432 670744
rect 3568 670704 364432 670732
rect 3568 670692 3574 670704
rect 364426 670692 364432 670704
rect 364484 670692 364490 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 362954 656928 362960 656940
rect 3476 656900 362960 656928
rect 3476 656888 3482 656900
rect 362954 656888 362960 656900
rect 363012 656888 363018 656940
rect 304994 643084 305000 643136
rect 305052 643124 305058 643136
rect 580166 643124 580172 643136
rect 305052 643096 580172 643124
rect 305052 643084 305058 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 367094 632108 367100 632120
rect 3476 632080 367100 632108
rect 3476 632068 3482 632080
rect 367094 632068 367100 632080
rect 367152 632068 367158 632120
rect 306374 630640 306380 630692
rect 306432 630680 306438 630692
rect 580166 630680 580172 630692
rect 306432 630652 580172 630680
rect 306432 630640 306438 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 369854 618304 369860 618316
rect 3200 618276 369860 618304
rect 3200 618264 3206 618276
rect 369854 618264 369860 618276
rect 369912 618264 369918 618316
rect 303614 616836 303620 616888
rect 303672 616876 303678 616888
rect 580166 616876 580172 616888
rect 303672 616848 580172 616876
rect 303672 616836 303678 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 368474 605860 368480 605872
rect 3292 605832 368480 605860
rect 3292 605820 3298 605832
rect 368474 605820 368480 605832
rect 368532 605820 368538 605872
rect 299566 590656 299572 590708
rect 299624 590696 299630 590708
rect 579798 590696 579804 590708
rect 299624 590668 579804 590696
rect 299624 590656 299630 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 372614 579680 372620 579692
rect 3384 579652 372620 579680
rect 3384 579640 3390 579652
rect 372614 579640 372620 579652
rect 372672 579640 372678 579692
rect 302234 576852 302240 576904
rect 302292 576892 302298 576904
rect 580166 576892 580172 576904
rect 302292 576864 580172 576892
rect 302292 576852 302298 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 375374 565876 375380 565888
rect 3476 565848 375380 565876
rect 3476 565836 3482 565848
rect 375374 565836 375380 565848
rect 375432 565836 375438 565888
rect 298094 563048 298100 563100
rect 298152 563088 298158 563100
rect 579798 563088 579804 563100
rect 298152 563060 579804 563088
rect 298152 563048 298158 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 373994 553432 374000 553444
rect 3476 553404 374000 553432
rect 3476 553392 3482 553404
rect 373994 553392 374000 553404
rect 374052 553392 374058 553444
rect 295334 536800 295340 536852
rect 295392 536840 295398 536852
rect 580166 536840 580172 536852
rect 295392 536812 580172 536840
rect 295392 536800 295398 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 376754 527184 376760 527196
rect 3476 527156 376760 527184
rect 3476 527144 3482 527156
rect 376754 527144 376760 527156
rect 376812 527144 376818 527196
rect 296714 524424 296720 524476
rect 296772 524464 296778 524476
rect 580166 524464 580172 524476
rect 296772 524436 580172 524464
rect 296772 524424 296778 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 380986 514808 380992 514820
rect 3476 514780 380992 514808
rect 3476 514768 3482 514780
rect 380986 514768 380992 514780
rect 381044 514768 381050 514820
rect 293310 510620 293316 510672
rect 293368 510660 293374 510672
rect 580166 510660 580172 510672
rect 293368 510632 580172 510660
rect 293368 510620 293374 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 276014 502392 276020 502444
rect 276072 502432 276078 502444
rect 579246 502432 579252 502444
rect 276072 502404 579252 502432
rect 276072 502392 276078 502404
rect 579246 502392 579252 502404
rect 579304 502392 579310 502444
rect 270494 502324 270500 502376
rect 270552 502364 270558 502376
rect 579154 502364 579160 502376
rect 270552 502336 579160 502364
rect 270552 502324 270558 502336
rect 579154 502324 579160 502336
rect 579212 502324 579218 502376
rect 330846 502188 330852 502240
rect 330904 502228 330910 502240
rect 364334 502228 364340 502240
rect 330904 502200 364340 502228
rect 330904 502188 330910 502200
rect 364334 502188 364340 502200
rect 364392 502188 364398 502240
rect 299474 502120 299480 502172
rect 299532 502160 299538 502172
rect 335538 502160 335544 502172
rect 299532 502132 335544 502160
rect 299532 502120 299538 502132
rect 335538 502120 335544 502132
rect 335596 502120 335602 502172
rect 325602 502052 325608 502104
rect 325660 502092 325666 502104
rect 429194 502092 429200 502104
rect 325660 502064 429200 502092
rect 325660 502052 325666 502064
rect 429194 502052 429200 502064
rect 429252 502052 429258 502104
rect 234614 501984 234620 502036
rect 234672 502024 234678 502036
rect 340874 502024 340880 502036
rect 234672 501996 340880 502024
rect 234672 501984 234678 501996
rect 340874 501984 340880 501996
rect 340932 501984 340938 502036
rect 322106 501916 322112 501968
rect 322164 501956 322170 501968
rect 462314 501956 462320 501968
rect 322164 501928 462320 501956
rect 322164 501916 322170 501928
rect 462314 501916 462320 501928
rect 462372 501916 462378 501968
rect 320082 501848 320088 501900
rect 320140 501888 320146 501900
rect 494054 501888 494060 501900
rect 320140 501860 494060 501888
rect 320140 501848 320146 501860
rect 494054 501848 494060 501860
rect 494112 501848 494118 501900
rect 169754 501780 169760 501832
rect 169812 501820 169818 501832
rect 346026 501820 346032 501832
rect 169812 501792 346032 501820
rect 169812 501780 169818 501792
rect 346026 501780 346032 501792
rect 346084 501780 346090 501832
rect 315114 501712 315120 501764
rect 315172 501752 315178 501764
rect 558914 501752 558920 501764
rect 315172 501724 558920 501752
rect 315172 501712 315178 501724
rect 558914 501712 558920 501724
rect 558972 501712 558978 501764
rect 104894 501644 104900 501696
rect 104952 501684 104958 501696
rect 351270 501684 351276 501696
rect 104952 501656 351276 501684
rect 104952 501644 104958 501656
rect 351270 501644 351276 501656
rect 351328 501644 351334 501696
rect 40034 501576 40040 501628
rect 40092 501616 40098 501628
rect 356514 501616 356520 501628
rect 40092 501588 356520 501616
rect 40092 501576 40098 501588
rect 356514 501576 356520 501588
rect 356572 501576 356578 501628
rect 265986 501168 265992 501220
rect 266044 501208 266050 501220
rect 579062 501208 579068 501220
rect 266044 501180 579068 501208
rect 266044 501168 266050 501180
rect 579062 501168 579068 501180
rect 579120 501168 579126 501220
rect 260558 501100 260564 501152
rect 260616 501140 260622 501152
rect 578970 501140 578976 501152
rect 260616 501112 578976 501140
rect 260616 501100 260622 501112
rect 578970 501100 578976 501112
rect 579028 501100 579034 501152
rect 255222 501032 255228 501084
rect 255280 501072 255286 501084
rect 578878 501072 578884 501084
rect 255280 501044 578884 501072
rect 255280 501032 255286 501044
rect 578878 501032 578884 501044
rect 578936 501032 578942 501084
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 358722 501004 358728 501016
rect 3108 500976 358728 501004
rect 3108 500964 3114 500976
rect 358722 500964 358728 500976
rect 358780 500964 358786 501016
rect 335998 500896 336004 500948
rect 336056 500936 336062 500948
rect 337286 500936 337292 500948
rect 336056 500908 337292 500936
rect 336056 500896 336062 500908
rect 337286 500896 337292 500908
rect 337344 500896 337350 500948
rect 337378 500896 337384 500948
rect 337436 500936 337442 500948
rect 342530 500936 342536 500948
rect 337436 500908 342536 500936
rect 337436 500896 337442 500908
rect 342530 500896 342536 500908
rect 342588 500896 342594 500948
rect 348418 500896 348424 500948
rect 348476 500936 348482 500948
rect 353294 500936 353300 500948
rect 348476 500908 353300 500936
rect 348476 500896 348482 500908
rect 353294 500896 353300 500908
rect 353352 500896 353358 500948
rect 355318 500896 355324 500948
rect 355376 500936 355382 500948
rect 360194 500936 360200 500948
rect 355376 500908 360200 500936
rect 355376 500896 355382 500908
rect 360194 500896 360200 500908
rect 360252 500896 360258 500948
rect 338758 500828 338764 500880
rect 338816 500868 338822 500880
rect 344278 500868 344284 500880
rect 338816 500840 344284 500868
rect 338816 500828 338822 500840
rect 344278 500828 344284 500840
rect 344336 500828 344342 500880
rect 353938 500488 353944 500540
rect 353996 500528 354002 500540
rect 358262 500528 358268 500540
rect 353996 500500 358268 500528
rect 353996 500488 354002 500500
rect 358262 500488 358268 500500
rect 358320 500488 358326 500540
rect 342898 500420 342904 500472
rect 342956 500460 342962 500472
rect 347958 500460 347964 500472
rect 342956 500432 347964 500460
rect 342956 500420 342962 500432
rect 347958 500420 347964 500432
rect 348016 500420 348022 500472
rect 349798 500420 349804 500472
rect 349856 500460 349862 500472
rect 354766 500460 354772 500472
rect 349856 500432 354772 500460
rect 349856 500420 349862 500432
rect 354766 500420 354772 500432
rect 354824 500420 354830 500472
rect 282914 500352 282920 500404
rect 282972 500392 282978 500404
rect 339034 500392 339040 500404
rect 282972 500364 339040 500392
rect 282972 500352 282978 500364
rect 339034 500352 339040 500364
rect 339092 500352 339098 500404
rect 344370 500352 344376 500404
rect 344428 500392 344434 500404
rect 349522 500392 349528 500404
rect 344428 500364 349528 500392
rect 344428 500352 344434 500364
rect 349522 500352 349528 500364
rect 349580 500352 349586 500404
rect 358722 500352 358728 500404
rect 358780 500392 358786 500404
rect 379514 500392 379520 500404
rect 358780 500364 379520 500392
rect 358780 500352 358786 500364
rect 379514 500352 379520 500364
rect 379572 500352 379578 500404
rect 234338 500284 234344 500336
rect 234396 500324 234402 500336
rect 409138 500324 409144 500336
rect 234396 500296 409144 500324
rect 234396 500284 234402 500296
rect 409138 500284 409144 500296
rect 409196 500284 409202 500336
rect 316862 500216 316868 500268
rect 316920 500256 316926 500268
rect 527174 500256 527180 500268
rect 316920 500228 527180 500256
rect 316920 500216 316926 500228
rect 527174 500216 527180 500228
rect 527232 500216 527238 500268
rect 267642 500148 267648 500200
rect 267700 500188 267706 500200
rect 578050 500188 578056 500200
rect 267700 500160 578056 500188
rect 267700 500148 267706 500160
rect 578050 500148 578056 500160
rect 578108 500148 578114 500200
rect 3234 500080 3240 500132
rect 3292 500120 3298 500132
rect 382826 500120 382832 500132
rect 3292 500092 382832 500120
rect 3292 500080 3298 500092
rect 382826 500080 382832 500092
rect 382884 500080 382890 500132
rect 4062 500012 4068 500064
rect 4120 500052 4126 500064
rect 384574 500052 384580 500064
rect 4120 500024 384580 500052
rect 4120 500012 4126 500024
rect 384574 500012 384580 500024
rect 384632 500012 384638 500064
rect 3326 499944 3332 499996
rect 3384 499984 3390 499996
rect 386598 499984 386604 499996
rect 3384 499956 386604 499984
rect 3384 499944 3390 499956
rect 386598 499944 386604 499956
rect 386656 499944 386662 499996
rect 3970 499876 3976 499928
rect 4028 499916 4034 499928
rect 388162 499916 388168 499928
rect 4028 499888 388168 499916
rect 4028 499876 4034 499888
rect 388162 499876 388168 499888
rect 388220 499876 388226 499928
rect 3786 499808 3792 499860
rect 3844 499848 3850 499860
rect 389910 499848 389916 499860
rect 3844 499820 389916 499848
rect 3844 499808 3850 499820
rect 389910 499808 389916 499820
rect 389968 499808 389974 499860
rect 3878 499740 3884 499792
rect 3936 499780 3942 499792
rect 391934 499780 391940 499792
rect 3936 499752 391940 499780
rect 3936 499740 3942 499752
rect 391934 499740 391940 499752
rect 391992 499740 391998 499792
rect 3694 499672 3700 499724
rect 3752 499712 3758 499724
rect 393406 499712 393412 499724
rect 3752 499684 393412 499712
rect 3752 499672 3758 499684
rect 393406 499672 393412 499684
rect 393464 499672 393470 499724
rect 3510 499604 3516 499656
rect 3568 499644 3574 499656
rect 395154 499644 395160 499656
rect 3568 499616 395160 499644
rect 3568 499604 3574 499616
rect 395154 499604 395160 499616
rect 395212 499604 395218 499656
rect 3602 499536 3608 499588
rect 3660 499576 3666 499588
rect 396902 499576 396908 499588
rect 3660 499548 396908 499576
rect 3660 499536 3666 499548
rect 396902 499536 396908 499548
rect 396960 499536 396966 499588
rect 233694 499060 233700 499112
rect 233752 499100 233758 499112
rect 402146 499100 402152 499112
rect 233752 499072 402152 499100
rect 233752 499060 233758 499072
rect 402146 499060 402152 499072
rect 402204 499060 402210 499112
rect 234430 498992 234436 499044
rect 234488 499032 234494 499044
rect 405734 499032 405740 499044
rect 234488 499004 405740 499032
rect 234488 498992 234494 499004
rect 405734 498992 405740 499004
rect 405792 498992 405798 499044
rect 234522 498924 234528 498976
rect 234580 498964 234586 498976
rect 407390 498964 407396 498976
rect 234580 498936 407396 498964
rect 234580 498924 234586 498936
rect 407390 498924 407396 498936
rect 407448 498924 407454 498976
rect 234154 498856 234160 498908
rect 234212 498896 234218 498908
rect 411254 498896 411260 498908
rect 234212 498868 411260 498896
rect 234212 498856 234218 498868
rect 411254 498856 411260 498868
rect 411312 498856 411318 498908
rect 234246 498788 234252 498840
rect 234304 498828 234310 498840
rect 412818 498828 412824 498840
rect 234304 498800 412824 498828
rect 234304 498788 234310 498800
rect 412818 498788 412824 498800
rect 412876 498788 412882 498840
rect 288802 498720 288808 498772
rect 288860 498760 288866 498772
rect 580902 498760 580908 498772
rect 288860 498732 580908 498760
rect 288860 498720 288866 498732
rect 580902 498720 580908 498732
rect 580960 498720 580966 498772
rect 274542 498652 274548 498704
rect 274600 498692 274606 498704
rect 577314 498692 577320 498704
rect 274600 498664 577320 498692
rect 274600 498652 274606 498664
rect 577314 498652 577320 498664
rect 577372 498652 577378 498704
rect 272978 498584 272984 498636
rect 273036 498624 273042 498636
rect 577406 498624 577412 498636
rect 273036 498596 577412 498624
rect 273036 498584 273042 498596
rect 577406 498584 577412 498596
rect 577464 498584 577470 498636
rect 269482 498516 269488 498568
rect 269540 498556 269546 498568
rect 578142 498556 578148 498568
rect 269540 498528 578148 498556
rect 269540 498516 269546 498528
rect 578142 498516 578148 498528
rect 578200 498516 578206 498568
rect 264238 498448 264244 498500
rect 264296 498488 264302 498500
rect 577958 498488 577964 498500
rect 264296 498460 577964 498488
rect 264296 498448 264302 498460
rect 577958 498448 577964 498460
rect 578016 498448 578022 498500
rect 258902 498380 258908 498432
rect 258960 498420 258966 498432
rect 577774 498420 577780 498432
rect 258960 498392 577780 498420
rect 258960 498380 258966 498392
rect 577774 498380 577780 498392
rect 577832 498380 577838 498432
rect 250162 498312 250168 498364
rect 250220 498352 250226 498364
rect 574830 498352 574836 498364
rect 250220 498324 574836 498352
rect 250220 498312 250226 498324
rect 574830 498312 574836 498324
rect 574888 498312 574894 498364
rect 253658 498244 253664 498296
rect 253716 498284 253722 498296
rect 577682 498284 577688 498296
rect 253716 498256 577688 498284
rect 253716 498244 253722 498256
rect 577682 498244 577688 498256
rect 577740 498244 577746 498296
rect 248092 498176 248098 498228
rect 248150 498216 248156 498228
rect 577498 498216 577504 498228
rect 248150 498188 577504 498216
rect 248150 498176 248156 498188
rect 577498 498176 577504 498188
rect 577556 498176 577562 498228
rect 278222 497428 278228 497480
rect 278280 497428 278286 497480
rect 279970 497428 279976 497480
rect 280028 497428 280034 497480
rect 281534 497428 281540 497480
rect 281592 497428 281598 497480
rect 283466 497428 283472 497480
rect 283524 497428 283530 497480
rect 285214 497428 285220 497480
rect 285272 497428 285278 497480
rect 286870 497428 286876 497480
rect 286928 497468 286934 497480
rect 286928 497440 287054 497468
rect 286928 497428 286934 497440
rect 278240 496856 278268 497428
rect 279988 496924 280016 497428
rect 281552 496992 281580 497428
rect 283484 497060 283512 497428
rect 285232 497128 285260 497428
rect 287026 497196 287054 497440
rect 290550 497428 290556 497480
rect 290608 497428 290614 497480
rect 292298 497428 292304 497480
rect 292356 497468 292362 497480
rect 292356 497440 296714 497468
rect 292356 497428 292362 497440
rect 290568 497264 290596 497428
rect 296686 497332 296714 497440
rect 580166 497332 580172 497344
rect 296686 497304 580172 497332
rect 580166 497292 580172 497304
rect 580224 497292 580230 497344
rect 580074 497264 580080 497276
rect 290568 497236 580080 497264
rect 580074 497224 580080 497236
rect 580132 497224 580138 497276
rect 580718 497196 580724 497208
rect 287026 497168 580724 497196
rect 580718 497156 580724 497168
rect 580776 497156 580782 497208
rect 580810 497128 580816 497140
rect 285232 497100 580816 497128
rect 580810 497088 580816 497100
rect 580868 497088 580874 497140
rect 580626 497060 580632 497072
rect 283484 497032 580632 497060
rect 580626 497020 580632 497032
rect 580684 497020 580690 497072
rect 580442 496992 580448 497004
rect 281552 496964 580448 496992
rect 580442 496952 580448 496964
rect 580500 496952 580506 497004
rect 580534 496924 580540 496936
rect 279988 496896 580540 496924
rect 580534 496884 580540 496896
rect 580592 496884 580598 496936
rect 580350 496856 580356 496868
rect 278240 496828 580356 496856
rect 580350 496816 580356 496828
rect 580408 496816 580414 496868
rect 235074 338240 235080 338292
rect 235132 338240 235138 338292
rect 235092 338020 235120 338240
rect 235074 337968 235080 338020
rect 235132 337968 235138 338020
rect 314700 337764 314706 337816
rect 314758 337804 314764 337816
rect 314930 337804 314936 337816
rect 314758 337776 314936 337804
rect 314758 337764 314764 337776
rect 314930 337764 314936 337776
rect 314988 337764 314994 337816
rect 259454 336744 259460 336796
rect 259512 336784 259518 336796
rect 259822 336784 259828 336796
rect 259512 336756 259828 336784
rect 259512 336744 259518 336756
rect 259822 336744 259828 336756
rect 259880 336744 259886 336796
rect 307938 336744 307944 336796
rect 307996 336784 308002 336796
rect 308122 336784 308128 336796
rect 307996 336756 308128 336784
rect 307996 336744 308002 336756
rect 308122 336744 308128 336756
rect 308180 336744 308186 336796
rect 321554 336744 321560 336796
rect 321612 336784 321618 336796
rect 321830 336784 321836 336796
rect 321612 336756 321836 336784
rect 321612 336744 321618 336756
rect 321830 336744 321836 336756
rect 321888 336744 321894 336796
rect 378060 336756 378640 336784
rect 173158 336676 173164 336728
rect 173216 336716 173222 336728
rect 270218 336716 270224 336728
rect 173216 336688 270224 336716
rect 173216 336676 173222 336688
rect 270218 336676 270224 336688
rect 270276 336676 270282 336728
rect 274634 336676 274640 336728
rect 274692 336716 274698 336728
rect 275094 336716 275100 336728
rect 274692 336688 275100 336716
rect 274692 336676 274698 336688
rect 275094 336676 275100 336688
rect 275152 336676 275158 336728
rect 304994 336676 305000 336728
rect 305052 336716 305058 336728
rect 339586 336716 339592 336728
rect 305052 336688 339592 336716
rect 305052 336676 305058 336688
rect 339586 336676 339592 336688
rect 339644 336676 339650 336728
rect 354674 336676 354680 336728
rect 354732 336716 354738 336728
rect 354950 336716 354956 336728
rect 354732 336688 354956 336716
rect 354732 336676 354738 336688
rect 354950 336676 354956 336688
rect 355008 336676 355014 336728
rect 360102 336676 360108 336728
rect 360160 336716 360166 336728
rect 360838 336716 360844 336728
rect 360160 336688 360844 336716
rect 360160 336676 360166 336688
rect 360838 336676 360844 336688
rect 360896 336676 360902 336728
rect 369762 336676 369768 336728
rect 369820 336716 369826 336728
rect 373258 336716 373264 336728
rect 369820 336688 373264 336716
rect 369820 336676 369826 336688
rect 373258 336676 373264 336688
rect 373316 336676 373322 336728
rect 373350 336676 373356 336728
rect 373408 336716 373414 336728
rect 378060 336716 378088 336756
rect 373408 336688 378088 336716
rect 373408 336676 373414 336688
rect 378134 336676 378140 336728
rect 378192 336716 378198 336728
rect 378502 336716 378508 336728
rect 378192 336688 378508 336716
rect 378192 336676 378198 336688
rect 378502 336676 378508 336688
rect 378560 336676 378566 336728
rect 378612 336716 378640 336756
rect 380250 336716 380256 336728
rect 378612 336688 380256 336716
rect 380250 336676 380256 336688
rect 380308 336676 380314 336728
rect 386322 336676 386328 336728
rect 386380 336716 386386 336728
rect 411898 336716 411904 336728
rect 386380 336688 411904 336716
rect 386380 336676 386386 336688
rect 411898 336676 411904 336688
rect 411956 336676 411962 336728
rect 414014 336676 414020 336728
rect 414072 336716 414078 336728
rect 414382 336716 414388 336728
rect 414072 336688 414388 336716
rect 414072 336676 414078 336688
rect 414382 336676 414388 336688
rect 414440 336676 414446 336728
rect 426434 336676 426440 336728
rect 426492 336716 426498 336728
rect 427170 336716 427176 336728
rect 426492 336688 427176 336716
rect 426492 336676 426498 336688
rect 427170 336676 427176 336688
rect 427228 336676 427234 336728
rect 428642 336676 428648 336728
rect 428700 336716 428706 336728
rect 451918 336716 451924 336728
rect 428700 336688 451924 336716
rect 428700 336676 428706 336688
rect 451918 336676 451924 336688
rect 451976 336676 451982 336728
rect 163498 336608 163504 336660
rect 163556 336648 163562 336660
rect 267826 336648 267832 336660
rect 163556 336620 267832 336648
rect 163556 336608 163562 336620
rect 267826 336608 267832 336620
rect 267884 336608 267890 336660
rect 298094 336608 298100 336660
rect 298152 336648 298158 336660
rect 337102 336648 337108 336660
rect 298152 336620 337108 336648
rect 298152 336608 298158 336620
rect 337102 336608 337108 336620
rect 337160 336608 337166 336660
rect 360010 336608 360016 336660
rect 360068 336648 360074 336660
rect 362954 336648 362960 336660
rect 360068 336620 362960 336648
rect 360068 336608 360074 336620
rect 362954 336608 362960 336620
rect 363012 336608 363018 336660
rect 373718 336608 373724 336660
rect 373776 336648 373782 336660
rect 400766 336648 400772 336660
rect 373776 336620 400772 336648
rect 373776 336608 373782 336620
rect 400766 336608 400772 336620
rect 400824 336608 400830 336660
rect 433518 336608 433524 336660
rect 433576 336648 433582 336660
rect 458818 336648 458824 336660
rect 433576 336620 458824 336648
rect 433576 336608 433582 336620
rect 458818 336608 458824 336620
rect 458876 336608 458882 336660
rect 153838 336540 153844 336592
rect 153896 336580 153902 336592
rect 265342 336580 265348 336592
rect 153896 336552 265348 336580
rect 153896 336540 153902 336552
rect 265342 336540 265348 336552
rect 265400 336540 265406 336592
rect 291194 336540 291200 336592
rect 291252 336580 291258 336592
rect 328914 336580 328920 336592
rect 291252 336552 328920 336580
rect 291252 336540 291258 336552
rect 328914 336540 328920 336552
rect 328972 336540 328978 336592
rect 333514 336580 333520 336592
rect 329024 336552 333520 336580
rect 149698 336472 149704 336524
rect 149756 336512 149762 336524
rect 264054 336512 264060 336524
rect 149756 336484 264060 336512
rect 149756 336472 149762 336484
rect 264054 336472 264060 336484
rect 264112 336472 264118 336524
rect 287054 336472 287060 336524
rect 287112 336512 287118 336524
rect 329024 336512 329052 336552
rect 333514 336540 333520 336552
rect 333572 336540 333578 336592
rect 345382 336540 345388 336592
rect 345440 336580 345446 336592
rect 353386 336580 353392 336592
rect 345440 336552 353392 336580
rect 345440 336540 345446 336552
rect 353386 336540 353392 336552
rect 353444 336540 353450 336592
rect 364978 336540 364984 336592
rect 365036 336580 365042 336592
rect 377398 336580 377404 336592
rect 365036 336552 377404 336580
rect 365036 336540 365042 336552
rect 377398 336540 377404 336552
rect 377456 336540 377462 336592
rect 388438 336540 388444 336592
rect 388496 336580 388502 336592
rect 416038 336580 416044 336592
rect 388496 336552 416044 336580
rect 388496 336540 388502 336552
rect 416038 336540 416044 336552
rect 416096 336540 416102 336592
rect 434622 336540 434628 336592
rect 434680 336580 434686 336592
rect 472618 336580 472624 336592
rect 434680 336552 472624 336580
rect 434680 336540 434686 336552
rect 472618 336540 472624 336552
rect 472676 336540 472682 336592
rect 332226 336512 332232 336524
rect 287112 336484 329052 336512
rect 329116 336484 332232 336512
rect 287112 336472 287118 336484
rect 145558 336404 145564 336456
rect 145616 336444 145622 336456
rect 261662 336444 261668 336456
rect 145616 336416 261668 336444
rect 145616 336404 145622 336416
rect 261662 336404 261668 336416
rect 261720 336404 261726 336456
rect 284294 336404 284300 336456
rect 284352 336444 284358 336456
rect 329116 336444 329144 336484
rect 332226 336472 332232 336484
rect 332284 336472 332290 336524
rect 366450 336472 366456 336524
rect 366508 336512 366514 336524
rect 379974 336512 379980 336524
rect 366508 336484 379980 336512
rect 366508 336472 366514 336484
rect 379974 336472 379980 336484
rect 380032 336472 380038 336524
rect 389726 336472 389732 336524
rect 389784 336512 389790 336524
rect 433978 336512 433984 336524
rect 389784 336484 433984 336512
rect 389784 336472 389790 336484
rect 433978 336472 433984 336484
rect 434036 336472 434042 336524
rect 284352 336416 329144 336444
rect 284352 336404 284358 336416
rect 331858 336404 331864 336456
rect 331916 336444 331922 336456
rect 345014 336444 345020 336456
rect 331916 336416 345020 336444
rect 331916 336404 331922 336416
rect 345014 336404 345020 336416
rect 345072 336404 345078 336456
rect 375282 336404 375288 336456
rect 375340 336444 375346 336456
rect 402238 336444 402244 336456
rect 375340 336416 402244 336444
rect 375340 336404 375346 336416
rect 402238 336404 402244 336416
rect 402296 336404 402302 336456
rect 426618 336404 426624 336456
rect 426676 336444 426682 336456
rect 475378 336444 475384 336456
rect 426676 336416 475384 336444
rect 426676 336404 426682 336416
rect 475378 336404 475384 336416
rect 475436 336404 475442 336456
rect 45554 336336 45560 336388
rect 45612 336376 45618 336388
rect 250714 336376 250720 336388
rect 45612 336348 250720 336376
rect 45612 336336 45618 336348
rect 250714 336336 250720 336348
rect 250772 336336 250778 336388
rect 262950 336336 262956 336388
rect 263008 336376 263014 336388
rect 315206 336376 315212 336388
rect 263008 336348 315212 336376
rect 263008 336336 263014 336348
rect 315206 336336 315212 336348
rect 315264 336336 315270 336388
rect 316034 336336 316040 336388
rect 316092 336376 316098 336388
rect 343174 336376 343180 336388
rect 316092 336348 343180 336376
rect 316092 336336 316098 336348
rect 343174 336336 343180 336348
rect 343232 336336 343238 336388
rect 368566 336336 368572 336388
rect 368624 336376 368630 336388
rect 384298 336376 384304 336388
rect 368624 336348 384304 336376
rect 368624 336336 368630 336348
rect 384298 336336 384304 336348
rect 384356 336336 384362 336388
rect 394602 336336 394608 336388
rect 394660 336376 394666 336388
rect 460198 336376 460204 336388
rect 394660 336348 460204 336376
rect 394660 336336 394666 336348
rect 460198 336336 460204 336348
rect 460256 336336 460262 336388
rect 38654 336268 38660 336320
rect 38712 336308 38718 336320
rect 248414 336308 248420 336320
rect 38712 336280 248420 336308
rect 38712 336268 38718 336280
rect 248414 336268 248420 336280
rect 248472 336268 248478 336320
rect 264238 336268 264244 336320
rect 264296 336308 264302 336320
rect 318886 336308 318892 336320
rect 264296 336280 318892 336308
rect 264296 336268 264302 336280
rect 318886 336268 318892 336280
rect 318944 336268 318950 336320
rect 328914 336268 328920 336320
rect 328972 336308 328978 336320
rect 334710 336308 334716 336320
rect 328972 336280 334716 336308
rect 328972 336268 328978 336280
rect 334710 336268 334716 336280
rect 334768 336268 334774 336320
rect 347314 336308 347320 336320
rect 334820 336280 347320 336308
rect 31754 336200 31760 336252
rect 31812 336240 31818 336252
rect 245838 336240 245844 336252
rect 31812 336212 245844 336240
rect 31812 336200 31818 336212
rect 245838 336200 245844 336212
rect 245896 336200 245902 336252
rect 273622 336200 273628 336252
rect 273680 336240 273686 336252
rect 328730 336240 328736 336252
rect 273680 336212 328736 336240
rect 273680 336200 273686 336212
rect 328730 336200 328736 336212
rect 328788 336200 328794 336252
rect 24854 336132 24860 336184
rect 24912 336172 24918 336184
rect 243446 336172 243452 336184
rect 24912 336144 243452 336172
rect 24912 336132 24918 336144
rect 243446 336132 243452 336144
rect 243504 336132 243510 336184
rect 261478 336132 261484 336184
rect 261536 336172 261542 336184
rect 319714 336172 319720 336184
rect 261536 336144 319720 336172
rect 261536 336132 261542 336144
rect 319714 336132 319720 336144
rect 319772 336132 319778 336184
rect 327350 336132 327356 336184
rect 327408 336172 327414 336184
rect 334820 336172 334848 336280
rect 347314 336268 347320 336280
rect 347372 336268 347378 336320
rect 369854 336268 369860 336320
rect 369912 336308 369918 336320
rect 388438 336308 388444 336320
rect 369912 336280 388444 336308
rect 369912 336268 369918 336280
rect 388438 336268 388444 336280
rect 388496 336268 388502 336320
rect 393314 336268 393320 336320
rect 393372 336308 393378 336320
rect 460934 336308 460940 336320
rect 393372 336280 460940 336308
rect 393372 336268 393378 336280
rect 460934 336268 460940 336280
rect 460992 336268 460998 336320
rect 334986 336200 334992 336252
rect 335044 336240 335050 336252
rect 347774 336240 347780 336252
rect 335044 336212 347780 336240
rect 335044 336200 335050 336212
rect 347774 336200 347780 336212
rect 347832 336200 347838 336252
rect 371050 336200 371056 336252
rect 371108 336240 371114 336252
rect 396074 336240 396080 336252
rect 371108 336212 396080 336240
rect 371108 336200 371114 336212
rect 396074 336200 396080 336212
rect 396132 336200 396138 336252
rect 399386 336200 399392 336252
rect 399444 336240 399450 336252
rect 468478 336240 468484 336252
rect 399444 336212 468484 336240
rect 399444 336200 399450 336212
rect 468478 336200 468484 336212
rect 468536 336200 468542 336252
rect 327408 336144 334848 336172
rect 327408 336132 327414 336144
rect 334894 336132 334900 336184
rect 334952 336172 334958 336184
rect 346854 336172 346860 336184
rect 334952 336144 346860 336172
rect 334952 336132 334958 336144
rect 346854 336132 346860 336144
rect 346912 336132 346918 336184
rect 372982 336132 372988 336184
rect 373040 336172 373046 336184
rect 393958 336172 393964 336184
rect 373040 336144 393964 336172
rect 373040 336132 373046 336144
rect 393958 336132 393964 336144
rect 394016 336132 394022 336184
rect 395982 336132 395988 336184
rect 396040 336172 396046 336184
rect 465718 336172 465724 336184
rect 396040 336144 465724 336172
rect 396040 336132 396046 336144
rect 465718 336132 465724 336144
rect 465776 336132 465782 336184
rect 15194 336064 15200 336116
rect 15252 336104 15258 336116
rect 240134 336104 240140 336116
rect 15252 336076 240140 336104
rect 15252 336064 15258 336076
rect 240134 336064 240140 336076
rect 240192 336064 240198 336116
rect 269114 336064 269120 336116
rect 269172 336104 269178 336116
rect 327442 336104 327448 336116
rect 269172 336076 327448 336104
rect 269172 336064 269178 336076
rect 327442 336064 327448 336076
rect 327500 336064 327506 336116
rect 334618 336064 334624 336116
rect 334676 336104 334682 336116
rect 349522 336104 349528 336116
rect 334676 336076 349528 336104
rect 334676 336064 334682 336076
rect 349522 336064 349528 336076
rect 349580 336064 349586 336116
rect 377950 336064 377956 336116
rect 378008 336104 378014 336116
rect 404998 336104 405004 336116
rect 378008 336076 405004 336104
rect 378008 336064 378014 336076
rect 404998 336064 405004 336076
rect 405056 336064 405062 336116
rect 416682 336064 416688 336116
rect 416740 336104 416746 336116
rect 528554 336104 528560 336116
rect 416740 336076 528560 336104
rect 416740 336064 416746 336076
rect 528554 336064 528560 336076
rect 528612 336064 528618 336116
rect 5534 335996 5540 336048
rect 5592 336036 5598 336048
rect 236914 336036 236920 336048
rect 5592 336008 236920 336036
rect 5592 335996 5598 336008
rect 236914 335996 236920 336008
rect 236972 335996 236978 336048
rect 266354 335996 266360 336048
rect 266412 336036 266418 336048
rect 326154 336036 326160 336048
rect 266412 336008 326160 336036
rect 266412 335996 266418 336008
rect 326154 335996 326160 336008
rect 326212 335996 326218 336048
rect 331214 335996 331220 336048
rect 331272 336036 331278 336048
rect 348510 336036 348516 336048
rect 331272 336008 348516 336036
rect 331272 335996 331278 336008
rect 348510 335996 348516 336008
rect 348568 335996 348574 336048
rect 366818 335996 366824 336048
rect 366876 336036 366882 336048
rect 374730 336036 374736 336048
rect 366876 336008 374736 336036
rect 366876 335996 366882 336008
rect 374730 335996 374736 336008
rect 374788 335996 374794 336048
rect 376570 335996 376576 336048
rect 376628 336036 376634 336048
rect 406562 336036 406568 336048
rect 376628 336008 406568 336036
rect 376628 335996 376634 336008
rect 406562 335996 406568 336008
rect 406620 335996 406626 336048
rect 418890 335996 418896 336048
rect 418948 336036 418954 336048
rect 535454 336036 535460 336048
rect 418948 336008 535460 336036
rect 418948 335996 418954 336008
rect 535454 335996 535460 336008
rect 535512 335996 535518 336048
rect 177298 335928 177304 335980
rect 177356 335968 177362 335980
rect 271414 335968 271420 335980
rect 177356 335940 271420 335968
rect 177356 335928 177362 335940
rect 271414 335928 271420 335940
rect 271472 335928 271478 335980
rect 307754 335928 307760 335980
rect 307812 335968 307818 335980
rect 340414 335968 340420 335980
rect 307812 335940 340420 335968
rect 307812 335928 307818 335940
rect 340414 335928 340420 335940
rect 340472 335928 340478 335980
rect 373902 335928 373908 335980
rect 373960 335968 373966 335980
rect 373960 335940 378824 335968
rect 373960 335928 373966 335940
rect 181438 335860 181444 335912
rect 181496 335900 181502 335912
rect 273806 335900 273812 335912
rect 181496 335872 273812 335900
rect 181496 335860 181502 335872
rect 273806 335860 273812 335872
rect 273864 335860 273870 335912
rect 311894 335860 311900 335912
rect 311952 335900 311958 335912
rect 342254 335900 342260 335912
rect 311952 335872 342260 335900
rect 311952 335860 311958 335872
rect 342254 335860 342260 335872
rect 342312 335860 342318 335912
rect 370958 335860 370964 335912
rect 371016 335900 371022 335912
rect 374638 335900 374644 335912
rect 371016 335872 374644 335900
rect 371016 335860 371022 335872
rect 374638 335860 374644 335872
rect 374696 335860 374702 335912
rect 378796 335900 378824 335940
rect 380066 335928 380072 335980
rect 380124 335968 380130 335980
rect 406378 335968 406384 335980
rect 380124 335940 406384 335968
rect 380124 335928 380130 335940
rect 406378 335928 406384 335940
rect 406436 335928 406442 335980
rect 426342 335928 426348 335980
rect 426400 335968 426406 335980
rect 447778 335968 447784 335980
rect 426400 335940 447784 335968
rect 426400 335928 426406 335940
rect 447778 335928 447784 335940
rect 447836 335928 447842 335980
rect 398098 335900 398104 335912
rect 378796 335872 398104 335900
rect 398098 335860 398104 335872
rect 398156 335860 398162 335912
rect 412818 335860 412824 335912
rect 412876 335900 412882 335912
rect 434070 335900 434076 335912
rect 412876 335872 434076 335900
rect 412876 335860 412882 335872
rect 434070 335860 434076 335872
rect 434128 335860 434134 335912
rect 188338 335792 188344 335844
rect 188396 335832 188402 335844
rect 276382 335832 276388 335844
rect 188396 335804 276388 335832
rect 188396 335792 188402 335804
rect 276382 335792 276388 335804
rect 276440 335792 276446 335844
rect 318794 335792 318800 335844
rect 318852 335832 318858 335844
rect 344462 335832 344468 335844
rect 318852 335804 344468 335832
rect 318852 335792 318858 335804
rect 344462 335792 344468 335804
rect 344520 335792 344526 335844
rect 362126 335792 362132 335844
rect 362184 335832 362190 335844
rect 363598 335832 363604 335844
rect 362184 335804 363604 335832
rect 362184 335792 362190 335804
rect 363598 335792 363604 335804
rect 363656 335792 363662 335844
rect 376662 335792 376668 335844
rect 376720 335832 376726 335844
rect 391198 335832 391204 335844
rect 376720 335804 391204 335832
rect 376720 335792 376726 335804
rect 391198 335792 391204 335804
rect 391256 335792 391262 335844
rect 421374 335792 421380 335844
rect 421432 335832 421438 335844
rect 440878 335832 440884 335844
rect 421432 335804 440884 335832
rect 421432 335792 421438 335804
rect 440878 335792 440884 335804
rect 440936 335792 440942 335844
rect 236638 335724 236644 335776
rect 236696 335764 236702 335776
rect 277578 335764 277584 335776
rect 236696 335736 277584 335764
rect 236696 335724 236702 335736
rect 277578 335724 277584 335736
rect 277636 335724 277642 335776
rect 326338 335724 326344 335776
rect 326396 335764 326402 335776
rect 338114 335764 338120 335776
rect 326396 335736 338120 335764
rect 326396 335724 326402 335736
rect 338114 335724 338120 335736
rect 338172 335724 338178 335776
rect 375466 335724 375472 335776
rect 375524 335764 375530 335776
rect 389818 335764 389824 335776
rect 375524 335736 389824 335764
rect 375524 335724 375530 335736
rect 389818 335724 389824 335736
rect 389876 335724 389882 335776
rect 431034 335724 431040 335776
rect 431092 335764 431098 335776
rect 450538 335764 450544 335776
rect 431092 335736 450544 335764
rect 431092 335724 431098 335736
rect 450538 335724 450544 335736
rect 450596 335724 450602 335776
rect 260098 335656 260104 335708
rect 260156 335696 260162 335708
rect 294966 335696 294972 335708
rect 260156 335668 294972 335696
rect 260156 335656 260162 335668
rect 294966 335656 294972 335668
rect 295024 335656 295030 335708
rect 325970 335656 325976 335708
rect 326028 335696 326034 335708
rect 334894 335696 334900 335708
rect 326028 335668 334900 335696
rect 326028 335656 326034 335668
rect 334894 335656 334900 335668
rect 334952 335656 334958 335708
rect 374270 335656 374276 335708
rect 374328 335696 374334 335708
rect 387150 335696 387156 335708
rect 374328 335668 387156 335696
rect 374328 335656 374334 335668
rect 387150 335656 387156 335668
rect 387208 335656 387214 335708
rect 423766 335656 423772 335708
rect 423824 335696 423830 335708
rect 440970 335696 440976 335708
rect 423824 335668 440976 335696
rect 423824 335656 423830 335668
rect 440970 335656 440976 335668
rect 441028 335656 441034 335708
rect 329098 335588 329104 335640
rect 329156 335628 329162 335640
rect 339126 335628 339132 335640
rect 329156 335600 339132 335628
rect 329156 335588 329162 335600
rect 339126 335588 339132 335600
rect 339184 335588 339190 335640
rect 333238 335520 333244 335572
rect 333296 335560 333302 335572
rect 334986 335560 334992 335572
rect 333296 335532 334992 335560
rect 333296 335520 333302 335532
rect 334986 335520 334992 335532
rect 335044 335520 335050 335572
rect 371878 335384 371884 335436
rect 371936 335424 371942 335436
rect 376018 335424 376024 335436
rect 371936 335396 376024 335424
rect 371936 335384 371942 335396
rect 376018 335384 376024 335396
rect 376076 335384 376082 335436
rect 353938 335316 353944 335368
rect 353996 335356 354002 335368
rect 356054 335356 356060 335368
rect 353996 335328 356060 335356
rect 353996 335316 354002 335328
rect 356054 335316 356060 335328
rect 356112 335316 356118 335368
rect 266630 330760 266636 330812
rect 266688 330800 266694 330812
rect 266906 330800 266912 330812
rect 266688 330772 266912 330800
rect 266688 330760 266694 330772
rect 266906 330760 266912 330772
rect 266964 330760 266970 330812
rect 291470 330760 291476 330812
rect 291528 330760 291534 330812
rect 292758 330760 292764 330812
rect 292816 330760 292822 330812
rect 301038 330760 301044 330812
rect 301096 330760 301102 330812
rect 320358 330760 320364 330812
rect 320416 330760 320422 330812
rect 291488 330608 291516 330760
rect 292776 330608 292804 330760
rect 301056 330608 301084 330760
rect 320376 330608 320404 330760
rect 291470 330556 291476 330608
rect 291528 330556 291534 330608
rect 292758 330556 292764 330608
rect 292816 330556 292822 330608
rect 301038 330556 301044 330608
rect 301096 330556 301102 330608
rect 320358 330556 320364 330608
rect 320416 330556 320422 330608
rect 234798 330488 234804 330540
rect 234856 330528 234862 330540
rect 235350 330528 235356 330540
rect 234856 330500 235356 330528
rect 234856 330488 234862 330500
rect 235350 330488 235356 330500
rect 235408 330488 235414 330540
rect 238754 330488 238760 330540
rect 238812 330528 238818 330540
rect 239766 330528 239772 330540
rect 238812 330500 239772 330528
rect 238812 330488 238818 330500
rect 239766 330488 239772 330500
rect 239824 330488 239830 330540
rect 240226 330488 240232 330540
rect 240284 330528 240290 330540
rect 240962 330528 240968 330540
rect 240284 330500 240968 330528
rect 240284 330488 240290 330500
rect 240962 330488 240968 330500
rect 241020 330488 241026 330540
rect 244274 330488 244280 330540
rect 244332 330528 244338 330540
rect 244642 330528 244648 330540
rect 244332 330500 244648 330528
rect 244332 330488 244338 330500
rect 244642 330488 244648 330500
rect 244700 330488 244706 330540
rect 245838 330488 245844 330540
rect 245896 330528 245902 330540
rect 246666 330528 246672 330540
rect 245896 330500 246672 330528
rect 245896 330488 245902 330500
rect 246666 330488 246672 330500
rect 246724 330488 246730 330540
rect 249886 330488 249892 330540
rect 249944 330528 249950 330540
rect 250346 330528 250352 330540
rect 249944 330500 250352 330528
rect 249944 330488 249950 330500
rect 250346 330488 250352 330500
rect 250404 330488 250410 330540
rect 252554 330488 252560 330540
rect 252612 330528 252618 330540
rect 253566 330528 253572 330540
rect 252612 330500 253572 330528
rect 252612 330488 252618 330500
rect 253566 330488 253572 330500
rect 253624 330488 253630 330540
rect 255498 330488 255504 330540
rect 255556 330528 255562 330540
rect 256418 330528 256424 330540
rect 255556 330500 256424 330528
rect 255556 330488 255562 330500
rect 256418 330488 256424 330500
rect 256476 330488 256482 330540
rect 256786 330488 256792 330540
rect 256844 330528 256850 330540
rect 257614 330528 257620 330540
rect 256844 330500 257620 330528
rect 256844 330488 256850 330500
rect 257614 330488 257620 330500
rect 257672 330488 257678 330540
rect 258166 330488 258172 330540
rect 258224 330528 258230 330540
rect 258810 330528 258816 330540
rect 258224 330500 258816 330528
rect 258224 330488 258230 330500
rect 258810 330488 258816 330500
rect 258868 330488 258874 330540
rect 259546 330488 259552 330540
rect 259604 330528 259610 330540
rect 260006 330528 260012 330540
rect 259604 330500 260012 330528
rect 259604 330488 259610 330500
rect 260006 330488 260012 330500
rect 260064 330488 260070 330540
rect 262214 330488 262220 330540
rect 262272 330528 262278 330540
rect 262858 330528 262864 330540
rect 262272 330500 262864 330528
rect 262272 330488 262278 330500
rect 262858 330488 262864 330500
rect 262916 330488 262922 330540
rect 267826 330488 267832 330540
rect 267884 330528 267890 330540
rect 268562 330528 268568 330540
rect 267884 330500 268568 330528
rect 267884 330488 267890 330500
rect 268562 330488 268568 330500
rect 268620 330488 268626 330540
rect 270586 330488 270592 330540
rect 270644 330528 270650 330540
rect 271046 330528 271052 330540
rect 270644 330500 271052 330528
rect 270644 330488 270650 330500
rect 271046 330488 271052 330500
rect 271104 330488 271110 330540
rect 271874 330488 271880 330540
rect 271932 330528 271938 330540
rect 272610 330528 272616 330540
rect 271932 330500 272616 330528
rect 271932 330488 271938 330500
rect 272610 330488 272616 330500
rect 272668 330488 272674 330540
rect 273530 330488 273536 330540
rect 273588 330528 273594 330540
rect 274266 330528 274272 330540
rect 273588 330500 274272 330528
rect 273588 330488 273594 330500
rect 274266 330488 274272 330500
rect 274324 330488 274330 330540
rect 276198 330488 276204 330540
rect 276256 330528 276262 330540
rect 276658 330528 276664 330540
rect 276256 330500 276664 330528
rect 276256 330488 276262 330500
rect 276658 330488 276664 330500
rect 276716 330488 276722 330540
rect 278774 330488 278780 330540
rect 278832 330528 278838 330540
rect 279142 330528 279148 330540
rect 278832 330500 279148 330528
rect 278832 330488 278838 330500
rect 279142 330488 279148 330500
rect 279200 330488 279206 330540
rect 280246 330488 280252 330540
rect 280304 330528 280310 330540
rect 280706 330528 280712 330540
rect 280304 330500 280712 330528
rect 280304 330488 280310 330500
rect 280706 330488 280712 330500
rect 280764 330488 280770 330540
rect 283006 330488 283012 330540
rect 283064 330528 283070 330540
rect 283558 330528 283564 330540
rect 283064 330500 283564 330528
rect 283064 330488 283070 330500
rect 283558 330488 283564 330500
rect 283616 330488 283622 330540
rect 284386 330488 284392 330540
rect 284444 330528 284450 330540
rect 284754 330528 284760 330540
rect 284444 330500 284760 330528
rect 284444 330488 284450 330500
rect 284754 330488 284760 330500
rect 284812 330488 284818 330540
rect 285766 330488 285772 330540
rect 285824 330528 285830 330540
rect 286042 330528 286048 330540
rect 285824 330500 286048 330528
rect 285824 330488 285830 330500
rect 286042 330488 286048 330500
rect 286100 330488 286106 330540
rect 287238 330488 287244 330540
rect 287296 330528 287302 330540
rect 287606 330528 287612 330540
rect 287296 330500 287612 330528
rect 287296 330488 287302 330500
rect 287606 330488 287612 330500
rect 287664 330488 287670 330540
rect 288434 330488 288440 330540
rect 288492 330528 288498 330540
rect 288894 330528 288900 330540
rect 288492 330500 288900 330528
rect 288492 330488 288498 330500
rect 288894 330488 288900 330500
rect 288952 330488 288958 330540
rect 289814 330488 289820 330540
rect 289872 330528 289878 330540
rect 290458 330528 290464 330540
rect 289872 330500 290464 330528
rect 289872 330488 289878 330500
rect 290458 330488 290464 330500
rect 290516 330488 290522 330540
rect 291378 330488 291384 330540
rect 291436 330528 291442 330540
rect 292114 330528 292120 330540
rect 291436 330500 292120 330528
rect 291436 330488 291442 330500
rect 292114 330488 292120 330500
rect 292172 330488 292178 330540
rect 292666 330488 292672 330540
rect 292724 330528 292730 330540
rect 293310 330528 293316 330540
rect 292724 330500 293316 330528
rect 292724 330488 292730 330500
rect 293310 330488 293316 330500
rect 293368 330488 293374 330540
rect 294046 330488 294052 330540
rect 294104 330528 294110 330540
rect 294506 330528 294512 330540
rect 294104 330500 294512 330528
rect 294104 330488 294110 330500
rect 294506 330488 294512 330500
rect 294564 330488 294570 330540
rect 296806 330488 296812 330540
rect 296864 330528 296870 330540
rect 297358 330528 297364 330540
rect 296864 330500 297364 330528
rect 296864 330488 296870 330500
rect 297358 330488 297364 330500
rect 297416 330488 297422 330540
rect 298186 330488 298192 330540
rect 298244 330528 298250 330540
rect 298554 330528 298560 330540
rect 298244 330500 298560 330528
rect 298244 330488 298250 330500
rect 298554 330488 298560 330500
rect 298612 330488 298618 330540
rect 299566 330488 299572 330540
rect 299624 330528 299630 330540
rect 300210 330528 300216 330540
rect 299624 330500 300216 330528
rect 299624 330488 299630 330500
rect 300210 330488 300216 330500
rect 300268 330488 300274 330540
rect 300946 330488 300952 330540
rect 301004 330528 301010 330540
rect 301406 330528 301412 330540
rect 301004 330500 301412 330528
rect 301004 330488 301010 330500
rect 301406 330488 301412 330500
rect 301464 330488 301470 330540
rect 311986 330488 311992 330540
rect 312044 330528 312050 330540
rect 312354 330528 312360 330540
rect 312044 330500 312360 330528
rect 312044 330488 312050 330500
rect 312354 330488 312360 330500
rect 312412 330488 312418 330540
rect 313366 330488 313372 330540
rect 313424 330528 313430 330540
rect 314010 330528 314016 330540
rect 313424 330500 314016 330528
rect 313424 330488 313430 330500
rect 314010 330488 314016 330500
rect 314068 330488 314074 330540
rect 314746 330488 314752 330540
rect 314804 330528 314810 330540
rect 315666 330528 315672 330540
rect 314804 330500 315672 330528
rect 314804 330488 314810 330500
rect 315666 330488 315672 330500
rect 315724 330488 315730 330540
rect 316218 330488 316224 330540
rect 316276 330528 316282 330540
rect 316862 330528 316868 330540
rect 316276 330500 316868 330528
rect 316276 330488 316282 330500
rect 316862 330488 316868 330500
rect 316920 330488 316926 330540
rect 317414 330488 317420 330540
rect 317472 330528 317478 330540
rect 318058 330528 318064 330540
rect 317472 330500 318064 330528
rect 317472 330488 317478 330500
rect 318058 330488 318064 330500
rect 318116 330488 318122 330540
rect 320266 330488 320272 330540
rect 320324 330528 320330 330540
rect 320910 330528 320916 330540
rect 320324 330500 320916 330528
rect 320324 330488 320330 330500
rect 320910 330488 320916 330500
rect 320968 330488 320974 330540
rect 321646 330488 321652 330540
rect 321704 330528 321710 330540
rect 322106 330528 322112 330540
rect 321704 330500 322112 330528
rect 321704 330488 321710 330500
rect 322106 330488 322112 330500
rect 322164 330488 322170 330540
rect 324314 330488 324320 330540
rect 324372 330528 324378 330540
rect 325326 330528 325332 330540
rect 324372 330500 325332 330528
rect 324372 330488 324378 330500
rect 325326 330488 325332 330500
rect 325384 330488 325390 330540
rect 327166 330488 327172 330540
rect 327224 330528 327230 330540
rect 327810 330528 327816 330540
rect 327224 330500 327816 330528
rect 327224 330488 327230 330500
rect 327810 330488 327816 330500
rect 327868 330488 327874 330540
rect 328546 330488 328552 330540
rect 328604 330528 328610 330540
rect 329466 330528 329472 330540
rect 328604 330500 329472 330528
rect 328604 330488 328610 330500
rect 329466 330488 329472 330500
rect 329524 330488 329530 330540
rect 340966 330488 340972 330540
rect 341024 330528 341030 330540
rect 341610 330528 341616 330540
rect 341024 330500 341616 330528
rect 341024 330488 341030 330500
rect 341610 330488 341616 330500
rect 341668 330488 341674 330540
rect 345290 330488 345296 330540
rect 345348 330528 345354 330540
rect 346026 330528 346032 330540
rect 345348 330500 346032 330528
rect 345348 330488 345354 330500
rect 346026 330488 346032 330500
rect 346084 330488 346090 330540
rect 349338 330488 349344 330540
rect 349396 330528 349402 330540
rect 349706 330528 349712 330540
rect 349396 330500 349712 330528
rect 349396 330488 349402 330500
rect 349706 330488 349712 330500
rect 349764 330488 349770 330540
rect 360286 330488 360292 330540
rect 360344 330528 360350 330540
rect 360654 330528 360660 330540
rect 360344 330500 360660 330528
rect 360344 330488 360350 330500
rect 360654 330488 360660 330500
rect 360712 330488 360718 330540
rect 363046 330488 363052 330540
rect 363104 330528 363110 330540
rect 363322 330528 363328 330540
rect 363104 330500 363328 330528
rect 363104 330488 363110 330500
rect 363322 330488 363328 330500
rect 363380 330488 363386 330540
rect 367186 330488 367192 330540
rect 367244 330528 367250 330540
rect 367922 330528 367928 330540
rect 367244 330500 367928 330528
rect 367244 330488 367250 330500
rect 367922 330488 367928 330500
rect 367980 330488 367986 330540
rect 379606 330488 379612 330540
rect 379664 330528 379670 330540
rect 380158 330528 380164 330540
rect 379664 330500 380164 330528
rect 379664 330488 379670 330500
rect 380158 330488 380164 330500
rect 380216 330488 380222 330540
rect 382458 330488 382464 330540
rect 382516 330528 382522 330540
rect 383010 330528 383016 330540
rect 382516 330500 383016 330528
rect 382516 330488 382522 330500
rect 383010 330488 383016 330500
rect 383068 330488 383074 330540
rect 383654 330488 383660 330540
rect 383712 330528 383718 330540
rect 384574 330528 384580 330540
rect 383712 330500 384580 330528
rect 383712 330488 383718 330500
rect 384574 330488 384580 330500
rect 384632 330488 384638 330540
rect 386506 330488 386512 330540
rect 386564 330528 386570 330540
rect 387426 330528 387432 330540
rect 386564 330500 387432 330528
rect 386564 330488 386570 330500
rect 387426 330488 387432 330500
rect 387484 330488 387490 330540
rect 410058 330488 410064 330540
rect 410116 330528 410122 330540
rect 410978 330528 410984 330540
rect 410116 330500 410984 330528
rect 410116 330488 410122 330500
rect 410978 330488 410984 330500
rect 411036 330488 411042 330540
rect 411254 330488 411260 330540
rect 411312 330528 411318 330540
rect 411806 330528 411812 330540
rect 411312 330500 411812 330528
rect 411312 330488 411318 330500
rect 411806 330488 411812 330500
rect 411864 330488 411870 330540
rect 414106 330488 414112 330540
rect 414164 330528 414170 330540
rect 414658 330528 414664 330540
rect 414164 330500 414664 330528
rect 414164 330488 414170 330500
rect 414658 330488 414664 330500
rect 414716 330488 414722 330540
rect 427814 330488 427820 330540
rect 427872 330528 427878 330540
rect 428826 330528 428832 330540
rect 427872 330500 428832 330528
rect 427872 330488 427878 330500
rect 428826 330488 428832 330500
rect 428884 330488 428890 330540
rect 429194 330488 429200 330540
rect 429252 330528 429258 330540
rect 430022 330528 430028 330540
rect 429252 330500 430028 330528
rect 429252 330488 429258 330500
rect 430022 330488 430028 330500
rect 430080 330488 430086 330540
rect 430574 330488 430580 330540
rect 430632 330528 430638 330540
rect 431218 330528 431224 330540
rect 430632 330500 431224 330528
rect 430632 330488 430638 330500
rect 431218 330488 431224 330500
rect 431276 330488 431282 330540
rect 234706 330420 234712 330472
rect 234764 330460 234770 330472
rect 235718 330460 235724 330472
rect 234764 330432 235724 330460
rect 234764 330420 234770 330432
rect 235718 330420 235724 330432
rect 235776 330420 235782 330472
rect 244366 330420 244372 330472
rect 244424 330460 244430 330472
rect 245010 330460 245016 330472
rect 244424 330432 245016 330460
rect 244424 330420 244430 330432
rect 245010 330420 245016 330432
rect 245068 330420 245074 330472
rect 255314 330420 255320 330472
rect 255372 330460 255378 330472
rect 255958 330460 255964 330472
rect 255372 330432 255964 330460
rect 255372 330420 255378 330432
rect 255958 330420 255964 330432
rect 256016 330420 256022 330472
rect 259638 330420 259644 330472
rect 259696 330460 259702 330472
rect 260466 330460 260472 330472
rect 259696 330432 260472 330460
rect 259696 330420 259702 330432
rect 260466 330420 260472 330432
rect 260524 330420 260530 330472
rect 262306 330420 262312 330472
rect 262364 330460 262370 330472
rect 263318 330460 263324 330472
rect 262364 330432 263324 330460
rect 262364 330420 262370 330432
rect 263318 330420 263324 330432
rect 263376 330420 263382 330472
rect 276106 330420 276112 330472
rect 276164 330460 276170 330472
rect 277118 330460 277124 330472
rect 276164 330432 277124 330460
rect 276164 330420 276170 330432
rect 277118 330420 277124 330432
rect 277176 330420 277182 330472
rect 280338 330420 280344 330472
rect 280396 330460 280402 330472
rect 281166 330460 281172 330472
rect 280396 330432 281172 330460
rect 280396 330420 280402 330432
rect 281166 330420 281172 330432
rect 281224 330420 281230 330472
rect 284478 330420 284484 330472
rect 284536 330460 284542 330472
rect 285214 330460 285220 330472
rect 284536 330432 285220 330460
rect 284536 330420 284542 330432
rect 285214 330420 285220 330432
rect 285272 330420 285278 330472
rect 287146 330420 287152 330472
rect 287204 330460 287210 330472
rect 288066 330460 288072 330472
rect 287204 330432 288072 330460
rect 287204 330420 287210 330432
rect 288066 330420 288072 330432
rect 288124 330420 288130 330472
rect 288526 330420 288532 330472
rect 288584 330460 288590 330472
rect 289262 330460 289268 330472
rect 288584 330432 289268 330460
rect 288584 330420 288590 330432
rect 289262 330420 289268 330432
rect 289320 330420 289326 330472
rect 298278 330420 298284 330472
rect 298336 330460 298342 330472
rect 299014 330460 299020 330472
rect 298336 330432 299020 330460
rect 298336 330420 298342 330432
rect 299014 330420 299020 330432
rect 299072 330420 299078 330472
rect 312078 330420 312084 330472
rect 312136 330460 312142 330472
rect 312814 330460 312820 330472
rect 312136 330432 312820 330460
rect 312136 330420 312142 330432
rect 312814 330420 312820 330432
rect 312872 330420 312878 330472
rect 317506 330420 317512 330472
rect 317564 330460 317570 330472
rect 318426 330460 318432 330472
rect 317564 330432 318432 330460
rect 317564 330420 317570 330432
rect 318426 330420 318432 330432
rect 318484 330420 318490 330472
rect 360194 330420 360200 330472
rect 360252 330460 360258 330472
rect 361114 330460 361120 330472
rect 360252 330432 361120 330460
rect 360252 330420 360258 330432
rect 361114 330420 361120 330432
rect 361172 330420 361178 330472
rect 379698 330420 379704 330472
rect 379756 330460 379762 330472
rect 380526 330460 380532 330472
rect 379756 330432 380532 330460
rect 379756 330420 379762 330432
rect 380526 330420 380532 330432
rect 380584 330420 380590 330472
rect 382274 330420 382280 330472
rect 382332 330460 382338 330472
rect 383378 330460 383384 330472
rect 382332 330432 383384 330460
rect 382332 330420 382338 330432
rect 383378 330420 383384 330432
rect 383436 330420 383442 330472
rect 409874 330420 409880 330472
rect 409932 330460 409938 330472
rect 410610 330460 410616 330472
rect 409932 330432 410616 330460
rect 409932 330420 409938 330432
rect 410610 330420 410616 330432
rect 410668 330420 410674 330472
rect 411346 330420 411352 330472
rect 411404 330460 411410 330472
rect 412174 330460 412180 330472
rect 411404 330432 412180 330460
rect 411404 330420 411410 330432
rect 412174 330420 412180 330432
rect 412232 330420 412238 330472
rect 414198 330420 414204 330472
rect 414256 330460 414262 330472
rect 415026 330460 415032 330472
rect 414256 330432 415032 330460
rect 414256 330420 414262 330432
rect 415026 330420 415032 330432
rect 415084 330420 415090 330472
rect 430666 330420 430672 330472
rect 430724 330460 430730 330472
rect 431678 330460 431684 330472
rect 430724 330432 431684 330460
rect 430724 330420 430730 330432
rect 431678 330420 431684 330432
rect 431736 330420 431742 330472
rect 349246 330216 349252 330268
rect 349304 330256 349310 330268
rect 350074 330256 350080 330268
rect 349304 330228 350080 330256
rect 349304 330216 349310 330228
rect 350074 330216 350080 330228
rect 350132 330216 350138 330268
rect 258074 330080 258080 330132
rect 258132 330120 258138 330132
rect 258442 330120 258448 330132
rect 258132 330092 258448 330120
rect 258132 330080 258138 330092
rect 258442 330080 258448 330092
rect 258500 330080 258506 330132
rect 299474 330080 299480 330132
rect 299532 330120 299538 330132
rect 299842 330120 299848 330132
rect 299532 330092 299848 330120
rect 299532 330080 299538 330092
rect 299842 330080 299848 330092
rect 299900 330080 299906 330132
rect 253934 329944 253940 329996
rect 253992 329984 253998 329996
rect 254762 329984 254768 329996
rect 253992 329956 254768 329984
rect 253992 329944 253998 329956
rect 254762 329944 254768 329956
rect 254820 329944 254826 329996
rect 295334 329944 295340 329996
rect 295392 329984 295398 329996
rect 296162 329984 296168 329996
rect 295392 329956 296168 329984
rect 295392 329944 295398 329956
rect 296162 329944 296168 329956
rect 296220 329944 296226 329996
rect 416866 329672 416872 329724
rect 416924 329712 416930 329724
rect 417878 329712 417884 329724
rect 416924 329684 417884 329712
rect 416924 329672 416930 329684
rect 417878 329672 417884 329684
rect 417936 329672 417942 329724
rect 387794 329536 387800 329588
rect 387852 329576 387858 329588
rect 388622 329576 388628 329588
rect 387852 329548 388628 329576
rect 387852 329536 387858 329548
rect 388622 329536 388628 329548
rect 388680 329536 388686 329588
rect 256694 329128 256700 329180
rect 256752 329168 256758 329180
rect 257246 329168 257252 329180
rect 256752 329140 257252 329168
rect 256752 329128 256758 329140
rect 257246 329128 257252 329140
rect 257304 329128 257310 329180
rect 313274 328720 313280 328772
rect 313332 328760 313338 328772
rect 313642 328760 313648 328772
rect 313332 328732 313648 328760
rect 313332 328720 313338 328732
rect 313642 328720 313648 328732
rect 313700 328720 313706 328772
rect 365714 328720 365720 328772
rect 365772 328760 365778 328772
rect 366910 328760 366916 328772
rect 365772 328732 366916 328760
rect 365772 328720 365778 328732
rect 366910 328720 366916 328732
rect 366968 328720 366974 328772
rect 283098 328448 283104 328500
rect 283156 328488 283162 328500
rect 284018 328488 284024 328500
rect 283156 328460 284024 328488
rect 283156 328448 283162 328460
rect 284018 328448 284024 328460
rect 284076 328448 284082 328500
rect 363046 328312 363052 328364
rect 363104 328352 363110 328364
rect 363874 328352 363880 328364
rect 363104 328324 363880 328352
rect 363104 328312 363110 328324
rect 363874 328312 363880 328324
rect 363932 328312 363938 328364
rect 289906 327904 289912 327956
rect 289964 327944 289970 327956
rect 290918 327944 290924 327956
rect 289964 327916 290924 327944
rect 289964 327904 289970 327916
rect 290918 327904 290924 327916
rect 290976 327904 290982 327956
rect 329834 327768 329840 327820
rect 329892 327808 329898 327820
rect 330202 327808 330208 327820
rect 329892 327780 330208 327808
rect 329892 327768 329898 327780
rect 330202 327768 330208 327780
rect 330260 327768 330266 327820
rect 260926 327496 260932 327548
rect 260984 327536 260990 327548
rect 261294 327536 261300 327548
rect 260984 327508 261300 327536
rect 260984 327496 260990 327508
rect 261294 327496 261300 327508
rect 261352 327496 261358 327548
rect 408494 327292 408500 327344
rect 408552 327332 408558 327344
rect 409322 327332 409328 327344
rect 408552 327304 409328 327332
rect 408552 327292 408558 327304
rect 409322 327292 409328 327304
rect 409380 327292 409386 327344
rect 296898 327224 296904 327276
rect 296956 327264 296962 327276
rect 297818 327264 297824 327276
rect 296956 327236 297824 327264
rect 296956 327224 296962 327236
rect 297818 327224 297824 327236
rect 297876 327224 297882 327276
rect 325786 326884 325792 326936
rect 325844 326924 325850 326936
rect 326614 326924 326620 326936
rect 325844 326896 326620 326924
rect 325844 326884 325850 326896
rect 326614 326884 326620 326896
rect 326672 326884 326678 326936
rect 285674 326816 285680 326868
rect 285732 326856 285738 326868
rect 286410 326856 286416 326868
rect 285732 326828 286416 326856
rect 285732 326816 285738 326828
rect 286410 326816 286416 326828
rect 286468 326816 286474 326868
rect 329926 326816 329932 326868
rect 329984 326856 329990 326868
rect 330662 326856 330668 326868
rect 329984 326828 330668 326856
rect 329984 326816 329990 326828
rect 330662 326816 330668 326828
rect 330720 326816 330726 326868
rect 419718 326816 419724 326868
rect 419776 326816 419782 326868
rect 280154 326680 280160 326732
rect 280212 326720 280218 326732
rect 280522 326720 280528 326732
rect 280212 326692 280528 326720
rect 280212 326680 280218 326692
rect 280522 326680 280528 326692
rect 280580 326680 280586 326732
rect 309134 326680 309140 326732
rect 309192 326720 309198 326732
rect 309410 326720 309416 326732
rect 309192 326692 309416 326720
rect 309192 326680 309198 326692
rect 309410 326680 309416 326692
rect 309468 326680 309474 326732
rect 419736 326664 419764 326816
rect 419718 326612 419724 326664
rect 419776 326612 419782 326664
rect 396350 326476 396356 326528
rect 396408 326516 396414 326528
rect 396534 326516 396540 326528
rect 396408 326488 396540 326516
rect 396408 326476 396414 326488
rect 396534 326476 396540 326488
rect 396592 326476 396598 326528
rect 303614 326408 303620 326460
rect 303672 326448 303678 326460
rect 304718 326448 304724 326460
rect 303672 326420 304724 326448
rect 303672 326408 303678 326420
rect 304718 326408 304724 326420
rect 304776 326408 304782 326460
rect 305270 326408 305276 326460
rect 305328 326448 305334 326460
rect 305454 326448 305460 326460
rect 305328 326420 305460 326448
rect 305328 326408 305334 326420
rect 305454 326408 305460 326420
rect 305512 326408 305518 326460
rect 306558 326408 306564 326460
rect 306616 326408 306622 326460
rect 307938 326408 307944 326460
rect 307996 326448 308002 326460
rect 308766 326448 308772 326460
rect 307996 326420 308772 326448
rect 307996 326408 308002 326420
rect 308766 326408 308772 326420
rect 308824 326408 308830 326460
rect 310606 326408 310612 326460
rect 310664 326448 310670 326460
rect 311618 326448 311624 326460
rect 310664 326420 311624 326448
rect 310664 326408 310670 326420
rect 311618 326408 311624 326420
rect 311676 326408 311682 326460
rect 335538 326408 335544 326460
rect 335596 326448 335602 326460
rect 335814 326448 335820 326460
rect 335596 326420 335820 326448
rect 335596 326408 335602 326420
rect 335814 326408 335820 326420
rect 335872 326408 335878 326460
rect 352006 326408 352012 326460
rect 352064 326448 352070 326460
rect 352926 326448 352932 326460
rect 352064 326420 352932 326448
rect 352064 326408 352070 326420
rect 352926 326408 352932 326420
rect 352984 326408 352990 326460
rect 397638 326408 397644 326460
rect 397696 326448 397702 326460
rect 398374 326448 398380 326460
rect 397696 326420 398380 326448
rect 397696 326408 397702 326420
rect 398374 326408 398380 326420
rect 398432 326408 398438 326460
rect 404538 326408 404544 326460
rect 404596 326448 404602 326460
rect 405274 326448 405280 326460
rect 404596 326420 405280 326448
rect 404596 326408 404602 326420
rect 405274 326408 405280 326420
rect 405332 326408 405338 326460
rect 303798 326340 303804 326392
rect 303856 326380 303862 326392
rect 304258 326380 304264 326392
rect 303856 326352 304264 326380
rect 303856 326340 303862 326352
rect 304258 326340 304264 326352
rect 304316 326340 304322 326392
rect 305086 326340 305092 326392
rect 305144 326380 305150 326392
rect 305914 326380 305920 326392
rect 305144 326352 305920 326380
rect 305144 326340 305150 326352
rect 305914 326340 305920 326352
rect 305972 326340 305978 326392
rect 306576 326256 306604 326408
rect 307846 326340 307852 326392
rect 307904 326380 307910 326392
rect 308306 326380 308312 326392
rect 307904 326352 308312 326380
rect 307904 326340 307910 326352
rect 308306 326340 308312 326352
rect 308364 326340 308370 326392
rect 309226 326340 309232 326392
rect 309284 326380 309290 326392
rect 309962 326380 309968 326392
rect 309284 326352 309968 326380
rect 309284 326340 309290 326352
rect 309962 326340 309968 326352
rect 310020 326340 310026 326392
rect 310514 326340 310520 326392
rect 310572 326380 310578 326392
rect 311158 326380 311164 326392
rect 310572 326352 311164 326380
rect 310572 326340 310578 326352
rect 311158 326340 311164 326352
rect 311216 326340 311222 326392
rect 332686 326340 332692 326392
rect 332744 326380 332750 326392
rect 333054 326380 333060 326392
rect 332744 326352 333060 326380
rect 332744 326340 332750 326352
rect 333054 326340 333060 326352
rect 333112 326340 333118 326392
rect 335354 326340 335360 326392
rect 335412 326380 335418 326392
rect 335906 326380 335912 326392
rect 335412 326352 335912 326380
rect 335412 326340 335418 326352
rect 335906 326340 335912 326352
rect 335964 326340 335970 326392
rect 338206 326340 338212 326392
rect 338264 326380 338270 326392
rect 338758 326380 338764 326392
rect 338264 326352 338764 326380
rect 338264 326340 338270 326352
rect 338758 326340 338764 326352
rect 338816 326340 338822 326392
rect 350534 326340 350540 326392
rect 350592 326380 350598 326392
rect 351362 326380 351368 326392
rect 350592 326352 351368 326380
rect 350592 326340 350598 326352
rect 351362 326340 351368 326352
rect 351420 326340 351426 326392
rect 351914 326340 351920 326392
rect 351972 326380 351978 326392
rect 352558 326380 352564 326392
rect 351972 326352 352564 326380
rect 351972 326340 351978 326352
rect 352558 326340 352564 326352
rect 352616 326340 352622 326392
rect 353478 326340 353484 326392
rect 353536 326380 353542 326392
rect 354214 326380 354220 326392
rect 353536 326352 354220 326380
rect 353536 326340 353542 326352
rect 354214 326340 354220 326352
rect 354272 326340 354278 326392
rect 354766 326340 354772 326392
rect 354824 326380 354830 326392
rect 355410 326380 355416 326392
rect 354824 326352 355416 326380
rect 354824 326340 354830 326352
rect 355410 326340 355416 326352
rect 355468 326340 355474 326392
rect 389358 326340 389364 326392
rect 389416 326380 389422 326392
rect 390278 326380 390284 326392
rect 389416 326352 390284 326380
rect 389416 326340 389422 326352
rect 390278 326340 390284 326352
rect 390336 326340 390342 326392
rect 394694 326340 394700 326392
rect 394752 326380 394758 326392
rect 395154 326380 395160 326392
rect 394752 326352 395160 326380
rect 394752 326340 394758 326352
rect 395154 326340 395160 326352
rect 395212 326340 395218 326392
rect 396166 326340 396172 326392
rect 396224 326380 396230 326392
rect 396810 326380 396816 326392
rect 396224 326352 396816 326380
rect 396224 326340 396230 326352
rect 396810 326340 396816 326352
rect 396868 326340 396874 326392
rect 397454 326340 397460 326392
rect 397512 326380 397518 326392
rect 398006 326380 398012 326392
rect 397512 326352 398012 326380
rect 397512 326340 397518 326352
rect 398006 326340 398012 326352
rect 398064 326340 398070 326392
rect 398834 326340 398840 326392
rect 398892 326380 398898 326392
rect 399570 326380 399576 326392
rect 398892 326352 399576 326380
rect 398892 326340 398898 326352
rect 399570 326340 399576 326352
rect 399628 326340 399634 326392
rect 400214 326340 400220 326392
rect 400272 326380 400278 326392
rect 401226 326380 401232 326392
rect 400272 326352 401232 326380
rect 400272 326340 400278 326352
rect 401226 326340 401232 326352
rect 401284 326340 401290 326392
rect 402974 326340 402980 326392
rect 403032 326380 403038 326392
rect 403710 326380 403716 326392
rect 403032 326352 403716 326380
rect 403032 326340 403038 326352
rect 403710 326340 403716 326352
rect 403768 326340 403774 326392
rect 404354 326340 404360 326392
rect 404412 326380 404418 326392
rect 404906 326380 404912 326392
rect 404412 326352 404912 326380
rect 404412 326340 404418 326352
rect 404906 326340 404912 326352
rect 404964 326340 404970 326392
rect 405918 326340 405924 326392
rect 405976 326380 405982 326392
rect 406470 326380 406476 326392
rect 405976 326352 406476 326380
rect 405976 326340 405982 326352
rect 406470 326340 406476 326352
rect 406528 326340 406534 326392
rect 407206 326340 407212 326392
rect 407264 326380 407270 326392
rect 408126 326380 408132 326392
rect 407264 326352 408132 326380
rect 407264 326340 407270 326352
rect 408126 326340 408132 326352
rect 408184 326340 408190 326392
rect 418154 326340 418160 326392
rect 418212 326380 418218 326392
rect 419074 326380 419080 326392
rect 418212 326352 419080 326380
rect 418212 326340 418218 326352
rect 419074 326340 419080 326352
rect 419132 326340 419138 326392
rect 419626 326340 419632 326392
rect 419684 326380 419690 326392
rect 420270 326380 420276 326392
rect 419684 326352 420276 326380
rect 419684 326340 419690 326352
rect 420270 326340 420276 326352
rect 420328 326340 420334 326392
rect 420914 326340 420920 326392
rect 420972 326380 420978 326392
rect 421558 326380 421564 326392
rect 420972 326352 421564 326380
rect 420972 326340 420978 326352
rect 421558 326340 421564 326352
rect 421616 326340 421622 326392
rect 422294 326340 422300 326392
rect 422352 326380 422358 326392
rect 423122 326380 423128 326392
rect 422352 326352 423128 326380
rect 422352 326340 422358 326352
rect 423122 326340 423128 326352
rect 423180 326340 423186 326392
rect 242986 326204 242992 326256
rect 243044 326244 243050 326256
rect 243814 326244 243820 326256
rect 243044 326216 243820 326244
rect 243044 326204 243050 326216
rect 243814 326204 243820 326216
rect 243872 326204 243878 326256
rect 306558 326204 306564 326256
rect 306616 326204 306622 326256
rect 335538 326204 335544 326256
rect 335596 326244 335602 326256
rect 336366 326244 336372 326256
rect 335596 326216 336372 326244
rect 335596 326204 335602 326216
rect 336366 326204 336372 326216
rect 336424 326204 336430 326256
rect 400398 326204 400404 326256
rect 400456 326244 400462 326256
rect 400582 326244 400588 326256
rect 400456 326216 400588 326244
rect 400456 326204 400462 326216
rect 400582 326204 400588 326216
rect 400640 326204 400646 326256
rect 401594 325728 401600 325780
rect 401652 325768 401658 325780
rect 402422 325768 402428 325780
rect 401652 325740 402428 325768
rect 401652 325728 401658 325740
rect 402422 325728 402428 325740
rect 402480 325728 402486 325780
rect 577314 325456 577320 325508
rect 577372 325496 577378 325508
rect 580442 325496 580448 325508
rect 577372 325468 580448 325496
rect 577372 325456 577378 325468
rect 580442 325456 580448 325468
rect 580500 325456 580506 325508
rect 390646 325320 390652 325372
rect 390704 325360 390710 325372
rect 391474 325360 391480 325372
rect 390704 325332 391480 325360
rect 390704 325320 390710 325332
rect 391474 325320 391480 325332
rect 391532 325320 391538 325372
rect 400306 324232 400312 324284
rect 400364 324272 400370 324284
rect 400858 324272 400864 324284
rect 400364 324244 400864 324272
rect 400364 324232 400370 324244
rect 400858 324232 400864 324244
rect 400916 324232 400922 324284
rect 306466 323552 306472 323604
rect 306524 323592 306530 323604
rect 306650 323592 306656 323604
rect 306524 323564 306656 323592
rect 306524 323552 306530 323564
rect 306650 323552 306656 323564
rect 306708 323552 306714 323604
rect 352098 323552 352104 323604
rect 352156 323592 352162 323604
rect 352282 323592 352288 323604
rect 352156 323564 352288 323592
rect 352156 323552 352162 323564
rect 352282 323552 352288 323564
rect 352340 323552 352346 323604
rect 422386 323552 422392 323604
rect 422444 323592 422450 323604
rect 422570 323592 422576 323604
rect 422444 323564 422576 323592
rect 422444 323552 422450 323564
rect 422570 323552 422576 323564
rect 422628 323552 422634 323604
rect 425054 323416 425060 323468
rect 425112 323456 425118 323468
rect 425606 323456 425612 323468
rect 425112 323428 425612 323456
rect 425112 323416 425118 323428
rect 425606 323416 425612 323428
rect 425664 323416 425670 323468
rect 390554 323008 390560 323060
rect 390612 323048 390618 323060
rect 391106 323048 391112 323060
rect 390612 323020 391112 323048
rect 390612 323008 390618 323020
rect 391106 323008 391112 323020
rect 391164 323008 391170 323060
rect 306374 322736 306380 322788
rect 306432 322776 306438 322788
rect 307110 322776 307116 322788
rect 306432 322748 307116 322776
rect 306432 322736 306438 322748
rect 307110 322736 307116 322748
rect 307168 322736 307174 322788
rect 389174 322464 389180 322516
rect 389232 322504 389238 322516
rect 389910 322504 389916 322516
rect 389232 322476 389916 322504
rect 389232 322464 389238 322476
rect 389910 322464 389916 322476
rect 389968 322464 389974 322516
rect 423674 322464 423680 322516
rect 423732 322504 423738 322516
rect 424778 322504 424784 322516
rect 423732 322476 424784 322504
rect 423732 322464 423738 322476
rect 424778 322464 424784 322476
rect 424836 322464 424842 322516
rect 423766 322056 423772 322108
rect 423824 322096 423830 322108
rect 424318 322096 424324 322108
rect 423824 322068 424324 322096
rect 423824 322056 423830 322068
rect 424318 322056 424324 322068
rect 424376 322056 424382 322108
rect 403066 321648 403072 321700
rect 403124 321688 403130 321700
rect 403250 321688 403256 321700
rect 403124 321660 403256 321688
rect 403124 321648 403130 321660
rect 403250 321648 403256 321660
rect 403308 321648 403314 321700
rect 419534 319200 419540 319252
rect 419592 319240 419598 319252
rect 419810 319240 419816 319252
rect 419592 319212 419816 319240
rect 419592 319200 419598 319212
rect 419810 319200 419816 319212
rect 419868 319200 419874 319252
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 233694 306320 233700 306332
rect 3568 306292 233700 306320
rect 3568 306280 3574 306292
rect 233694 306280 233700 306292
rect 233752 306280 233758 306332
rect 577406 299412 577412 299464
rect 577464 299452 577470 299464
rect 579614 299452 579620 299464
rect 577464 299424 579620 299452
rect 577464 299412 577470 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 233786 293944 233792 293956
rect 3108 293916 233792 293944
rect 3108 293904 3114 293916
rect 233786 293904 233792 293916
rect 233844 293904 233850 293956
rect 578142 273164 578148 273216
rect 578200 273204 578206 273216
rect 579890 273204 579896 273216
rect 578200 273176 579896 273204
rect 578200 273164 578206 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 234522 255252 234528 255264
rect 3200 255224 234528 255252
rect 3200 255212 3206 255224
rect 234522 255212 234528 255224
rect 234580 255212 234586 255264
rect 578050 245556 578056 245608
rect 578108 245596 578114 245608
rect 579614 245596 579620 245608
rect 578108 245568 579620 245596
rect 578108 245556 578114 245568
rect 579614 245556 579620 245568
rect 579672 245556 579678 245608
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 234430 241448 234436 241460
rect 3568 241420 234436 241448
rect 3568 241408 3574 241420
rect 234430 241408 234436 241420
rect 234488 241408 234494 241460
rect 577958 233180 577964 233232
rect 578016 233220 578022 233232
rect 579798 233220 579804 233232
rect 578016 233192 579804 233220
rect 578016 233180 578022 233192
rect 579798 233180 579804 233192
rect 579856 233180 579862 233232
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 234338 215268 234344 215280
rect 3384 215240 234344 215268
rect 3384 215228 3390 215240
rect 234338 215228 234344 215240
rect 234396 215228 234402 215280
rect 577866 206932 577872 206984
rect 577924 206972 577930 206984
rect 579982 206972 579988 206984
rect 577924 206944 579988 206972
rect 577924 206932 577930 206944
rect 579982 206932 579988 206944
rect 580040 206932 580046 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 234246 202824 234252 202836
rect 3108 202796 234252 202824
rect 3108 202784 3114 202796
rect 234246 202784 234252 202796
rect 234304 202784 234310 202836
rect 577774 193128 577780 193180
rect 577832 193168 577838 193180
rect 579614 193168 579620 193180
rect 577832 193140 579620 193168
rect 577832 193128 577838 193140
rect 579614 193128 579620 193140
rect 579672 193128 579678 193180
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 234154 189020 234160 189032
rect 3568 188992 234160 189020
rect 3568 188980 3574 188992
rect 234154 188980 234160 188992
rect 234212 188980 234218 189032
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 234062 164200 234068 164212
rect 3292 164172 234068 164200
rect 3292 164160 3298 164172
rect 234062 164160 234068 164172
rect 234120 164160 234126 164212
rect 577682 153144 577688 153196
rect 577740 153184 577746 153196
rect 580626 153184 580632 153196
rect 577740 153156 580632 153184
rect 577740 153144 577746 153156
rect 580626 153144 580632 153156
rect 580684 153144 580690 153196
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 235074 150396 235080 150408
rect 3568 150368 235080 150396
rect 3568 150356 3574 150368
rect 235074 150356 235080 150368
rect 235132 150356 235138 150408
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 233970 137952 233976 137964
rect 3568 137924 233976 137952
rect 3568 137912 3574 137924
rect 233970 137912 233976 137924
rect 234028 137912 234034 137964
rect 577498 112956 577504 113008
rect 577556 112996 577562 113008
rect 580350 112996 580356 113008
rect 577556 112968 580356 112996
rect 577556 112956 577562 112968
rect 580350 112956 580356 112968
rect 580408 112956 580414 113008
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 233878 111772 233884 111784
rect 3200 111744 233884 111772
rect 3200 111732 3206 111744
rect 233878 111732 233884 111744
rect 233936 111732 233942 111784
rect 574830 100648 574836 100700
rect 574888 100688 574894 100700
rect 580166 100688 580172 100700
rect 574888 100660 580172 100688
rect 574888 100648 574894 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 577590 73108 577596 73160
rect 577648 73148 577654 73160
rect 579706 73148 579712 73160
rect 577648 73120 579712 73148
rect 577648 73108 577654 73120
rect 579706 73108 579712 73120
rect 579764 73108 579770 73160
rect 574738 60664 574744 60716
rect 574796 60704 574802 60716
rect 580166 60704 580172 60716
rect 574796 60676 580172 60704
rect 574796 60664 574802 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 74534 20204 74540 20256
rect 74592 20244 74598 20256
rect 259638 20244 259644 20256
rect 74592 20216 259644 20244
rect 74592 20204 74598 20216
rect 259638 20204 259644 20216
rect 259696 20204 259702 20256
rect 70394 20136 70400 20188
rect 70452 20176 70458 20188
rect 259730 20176 259736 20188
rect 70452 20148 259736 20176
rect 70452 20136 70458 20148
rect 259730 20136 259736 20148
rect 259788 20136 259794 20188
rect 67634 20068 67640 20120
rect 67692 20108 67698 20120
rect 258258 20108 258264 20120
rect 67692 20080 258264 20108
rect 67692 20068 67698 20080
rect 258258 20068 258264 20080
rect 258316 20068 258322 20120
rect 63494 20000 63500 20052
rect 63552 20040 63558 20052
rect 256878 20040 256884 20052
rect 63552 20012 256884 20040
rect 63552 20000 63558 20012
rect 256878 20000 256884 20012
rect 256936 20000 256942 20052
rect 60734 19932 60740 19984
rect 60792 19972 60798 19984
rect 255590 19972 255596 19984
rect 60792 19944 255596 19972
rect 60792 19932 60798 19944
rect 255590 19932 255596 19944
rect 255648 19932 255654 19984
rect 187694 19252 187700 19304
rect 187752 19292 187758 19304
rect 299658 19292 299664 19304
rect 187752 19264 299664 19292
rect 187752 19252 187758 19264
rect 299658 19252 299664 19264
rect 299716 19252 299722 19304
rect 151814 19184 151820 19236
rect 151872 19224 151878 19236
rect 287422 19224 287428 19236
rect 151872 19196 287428 19224
rect 151872 19184 151878 19196
rect 287422 19184 287428 19196
rect 287480 19184 287486 19236
rect 121454 19116 121460 19168
rect 121512 19156 121518 19168
rect 276198 19156 276204 19168
rect 121512 19128 276204 19156
rect 121512 19116 121518 19128
rect 276198 19116 276204 19128
rect 276256 19116 276262 19168
rect 118694 19048 118700 19100
rect 118752 19088 118758 19100
rect 274818 19088 274824 19100
rect 118752 19060 274824 19088
rect 118752 19048 118758 19060
rect 274818 19048 274824 19060
rect 274876 19048 274882 19100
rect 114554 18980 114560 19032
rect 114612 19020 114618 19032
rect 273530 19020 273536 19032
rect 114612 18992 273536 19020
rect 114612 18980 114618 18992
rect 273530 18980 273536 18992
rect 273588 18980 273594 19032
rect 56594 18912 56600 18964
rect 56652 18952 56658 18964
rect 254118 18952 254124 18964
rect 56652 18924 254124 18952
rect 56652 18912 56658 18924
rect 254118 18912 254124 18924
rect 254176 18912 254182 18964
rect 52454 18844 52460 18896
rect 52512 18884 52518 18896
rect 252830 18884 252836 18896
rect 52512 18856 252836 18884
rect 52512 18844 52518 18856
rect 252830 18844 252836 18856
rect 252888 18844 252894 18896
rect 49694 18776 49700 18828
rect 49752 18816 49758 18828
rect 251358 18816 251364 18828
rect 49752 18788 251364 18816
rect 49752 18776 49758 18788
rect 251358 18776 251364 18788
rect 251416 18776 251422 18828
rect 44174 18708 44180 18760
rect 44232 18748 44238 18760
rect 249886 18748 249892 18760
rect 44232 18720 249892 18748
rect 44232 18708 44238 18720
rect 249886 18708 249892 18720
rect 249944 18708 249950 18760
rect 41414 18640 41420 18692
rect 41472 18680 41478 18692
rect 248598 18680 248604 18692
rect 41472 18652 248604 18680
rect 41472 18640 41478 18652
rect 248598 18640 248604 18652
rect 248656 18640 248662 18692
rect 37274 18572 37280 18624
rect 37332 18612 37338 18624
rect 247218 18612 247224 18624
rect 37332 18584 247224 18612
rect 37332 18572 37338 18584
rect 247218 18572 247224 18584
rect 247276 18572 247282 18624
rect 191834 18504 191840 18556
rect 191892 18544 191898 18556
rect 301038 18544 301044 18556
rect 191892 18516 301044 18544
rect 191892 18504 191898 18516
rect 301038 18504 301044 18516
rect 301096 18504 301102 18556
rect 194594 18436 194600 18488
rect 194652 18476 194658 18488
rect 301130 18476 301136 18488
rect 194652 18448 301136 18476
rect 194652 18436 194658 18448
rect 301130 18436 301136 18448
rect 301188 18436 301194 18488
rect 198734 18368 198740 18420
rect 198792 18408 198798 18420
rect 302418 18408 302424 18420
rect 198792 18380 302424 18408
rect 198792 18368 198798 18380
rect 302418 18368 302424 18380
rect 302476 18368 302482 18420
rect 208394 17892 208400 17944
rect 208452 17932 208458 17944
rect 306558 17932 306564 17944
rect 208452 17904 306564 17932
rect 208452 17892 208458 17904
rect 306558 17892 306564 17904
rect 306616 17892 306622 17944
rect 204254 17824 204260 17876
rect 204312 17864 204318 17876
rect 305270 17864 305276 17876
rect 204312 17836 305276 17864
rect 204312 17824 204318 17836
rect 305270 17824 305276 17836
rect 305328 17824 305334 17876
rect 201494 17756 201500 17808
rect 201552 17796 201558 17808
rect 303890 17796 303896 17808
rect 201552 17768 303896 17796
rect 201552 17756 201558 17768
rect 303890 17756 303896 17768
rect 303948 17756 303954 17808
rect 197354 17688 197360 17740
rect 197412 17728 197418 17740
rect 302326 17728 302332 17740
rect 197412 17700 302332 17728
rect 197412 17688 197418 17700
rect 302326 17688 302332 17700
rect 302384 17688 302390 17740
rect 153194 17620 153200 17672
rect 153252 17660 153258 17672
rect 287238 17660 287244 17672
rect 153252 17632 287244 17660
rect 153252 17620 153258 17632
rect 287238 17620 287244 17632
rect 287296 17620 287302 17672
rect 150434 17552 150440 17604
rect 150492 17592 150498 17604
rect 285674 17592 285680 17604
rect 150492 17564 285680 17592
rect 150492 17552 150498 17564
rect 285674 17552 285680 17564
rect 285732 17552 285738 17604
rect 151906 17484 151912 17536
rect 151964 17524 151970 17536
rect 287330 17524 287336 17536
rect 151964 17496 287336 17524
rect 151964 17484 151970 17496
rect 287330 17484 287336 17496
rect 287388 17484 287394 17536
rect 149054 17416 149060 17468
rect 149112 17456 149118 17468
rect 285766 17456 285772 17468
rect 149112 17428 285772 17456
rect 149112 17416 149118 17428
rect 285766 17416 285772 17428
rect 285824 17416 285830 17468
rect 146294 17348 146300 17400
rect 146352 17388 146358 17400
rect 284478 17388 284484 17400
rect 146352 17360 284484 17388
rect 146352 17348 146358 17360
rect 284478 17348 284484 17360
rect 284536 17348 284542 17400
rect 147674 17280 147680 17332
rect 147732 17320 147738 17332
rect 285858 17320 285864 17332
rect 147732 17292 285864 17320
rect 147732 17280 147738 17292
rect 285858 17280 285864 17292
rect 285916 17280 285922 17332
rect 143534 17212 143540 17264
rect 143592 17252 143598 17264
rect 284570 17252 284576 17264
rect 143592 17224 284576 17252
rect 143592 17212 143598 17224
rect 284570 17212 284576 17224
rect 284628 17212 284634 17264
rect 211154 17144 211160 17196
rect 211212 17184 211218 17196
rect 308122 17184 308128 17196
rect 211212 17156 308128 17184
rect 211212 17144 211218 17156
rect 308122 17144 308128 17156
rect 308180 17144 308186 17196
rect 224954 17076 224960 17128
rect 225012 17116 225018 17128
rect 312170 17116 312176 17128
rect 225012 17088 312176 17116
rect 225012 17076 225018 17088
rect 312170 17076 312176 17088
rect 312228 17076 312234 17128
rect 227714 17008 227720 17060
rect 227772 17048 227778 17060
rect 313458 17048 313464 17060
rect 227772 17020 313464 17048
rect 227772 17008 227778 17020
rect 313458 17008 313464 17020
rect 313516 17008 313522 17060
rect 164418 16532 164424 16584
rect 164476 16572 164482 16584
rect 291470 16572 291476 16584
rect 164476 16544 291476 16572
rect 164476 16532 164482 16544
rect 291470 16532 291476 16544
rect 291528 16532 291534 16584
rect 161290 16464 161296 16516
rect 161348 16504 161354 16516
rect 290090 16504 290096 16516
rect 161348 16476 290096 16504
rect 161348 16464 161354 16476
rect 290090 16464 290096 16476
rect 290148 16464 290154 16516
rect 143626 16396 143632 16448
rect 143684 16436 143690 16448
rect 283098 16436 283104 16448
rect 143684 16408 283104 16436
rect 143684 16396 143690 16408
rect 283098 16396 283104 16408
rect 283156 16396 283162 16448
rect 125594 16328 125600 16380
rect 125652 16368 125658 16380
rect 277486 16368 277492 16380
rect 125652 16340 277492 16368
rect 125652 16328 125658 16340
rect 277486 16328 277492 16340
rect 277544 16328 277550 16380
rect 123018 16260 123024 16312
rect 123076 16300 123082 16312
rect 276106 16300 276112 16312
rect 123076 16272 276112 16300
rect 123076 16260 123082 16272
rect 276106 16260 276112 16272
rect 276164 16260 276170 16312
rect 119890 16192 119896 16244
rect 119948 16232 119954 16244
rect 276290 16232 276296 16244
rect 119948 16204 276296 16232
rect 119948 16192 119954 16204
rect 276290 16192 276296 16204
rect 276348 16192 276354 16244
rect 116394 16124 116400 16176
rect 116452 16164 116458 16176
rect 274726 16164 274732 16176
rect 116452 16136 274732 16164
rect 116452 16124 116458 16136
rect 274726 16124 274732 16136
rect 274784 16124 274790 16176
rect 112346 16056 112352 16108
rect 112404 16096 112410 16108
rect 273438 16096 273444 16108
rect 112404 16068 273444 16096
rect 112404 16056 112410 16068
rect 273438 16056 273444 16068
rect 273496 16056 273502 16108
rect 34514 15988 34520 16040
rect 34572 16028 34578 16040
rect 245838 16028 245844 16040
rect 34572 16000 245844 16028
rect 34572 15988 34578 16000
rect 245838 15988 245844 16000
rect 245896 15988 245902 16040
rect 30834 15920 30840 15972
rect 30892 15960 30898 15972
rect 245746 15960 245752 15972
rect 30892 15932 245752 15960
rect 30892 15920 30898 15932
rect 245746 15920 245752 15932
rect 245804 15920 245810 15972
rect 27706 15852 27712 15904
rect 27764 15892 27770 15904
rect 244458 15892 244464 15904
rect 27764 15864 244464 15892
rect 27764 15852 27770 15864
rect 244458 15852 244464 15864
rect 244516 15852 244522 15904
rect 168374 15784 168380 15836
rect 168432 15824 168438 15836
rect 292758 15824 292764 15836
rect 168432 15796 292764 15824
rect 168432 15784 168438 15796
rect 292758 15784 292764 15796
rect 292816 15784 292822 15836
rect 171962 15716 171968 15768
rect 172020 15756 172026 15768
rect 294138 15756 294144 15768
rect 172020 15728 294144 15756
rect 172020 15716 172026 15728
rect 294138 15716 294144 15728
rect 294196 15716 294202 15768
rect 221090 15648 221096 15700
rect 221148 15688 221154 15700
rect 310790 15688 310796 15700
rect 221148 15660 310796 15688
rect 221148 15648 221154 15660
rect 310790 15648 310796 15660
rect 310848 15648 310854 15700
rect 98178 15104 98184 15156
rect 98236 15144 98242 15156
rect 267826 15144 267832 15156
rect 98236 15116 267832 15144
rect 98236 15104 98242 15116
rect 267826 15104 267832 15116
rect 267884 15104 267890 15156
rect 93854 15036 93860 15088
rect 93912 15076 93918 15088
rect 266722 15076 266728 15088
rect 93912 15048 266728 15076
rect 93912 15036 93918 15048
rect 266722 15036 266728 15048
rect 266780 15036 266786 15088
rect 91554 14968 91560 15020
rect 91612 15008 91618 15020
rect 266630 15008 266636 15020
rect 91612 14980 266636 15008
rect 91612 14968 91618 14980
rect 266630 14968 266636 14980
rect 266688 14968 266694 15020
rect 87506 14900 87512 14952
rect 87564 14940 87570 14952
rect 265066 14940 265072 14952
rect 87564 14912 265072 14940
rect 87564 14900 87570 14912
rect 265066 14900 265072 14912
rect 265124 14900 265130 14952
rect 84194 14832 84200 14884
rect 84252 14872 84258 14884
rect 263686 14872 263692 14884
rect 84252 14844 263692 14872
rect 84252 14832 84258 14844
rect 263686 14832 263692 14844
rect 263744 14832 263750 14884
rect 80882 14764 80888 14816
rect 80940 14804 80946 14816
rect 262490 14804 262496 14816
rect 80940 14776 262496 14804
rect 80940 14764 80946 14776
rect 262490 14764 262496 14776
rect 262548 14764 262554 14816
rect 77386 14696 77392 14748
rect 77444 14736 77450 14748
rect 260926 14736 260932 14748
rect 77444 14708 260932 14736
rect 77444 14696 77450 14708
rect 260926 14696 260932 14708
rect 260984 14696 260990 14748
rect 73338 14628 73344 14680
rect 73396 14668 73402 14680
rect 259546 14668 259552 14680
rect 73396 14640 259552 14668
rect 73396 14628 73402 14640
rect 259546 14628 259552 14640
rect 259604 14628 259610 14680
rect 69842 14560 69848 14612
rect 69900 14600 69906 14612
rect 258166 14600 258172 14612
rect 69900 14572 258172 14600
rect 69900 14560 69906 14572
rect 258166 14560 258172 14572
rect 258224 14560 258230 14612
rect 66714 14492 66720 14544
rect 66772 14532 66778 14544
rect 256786 14532 256792 14544
rect 66772 14504 256792 14532
rect 66772 14492 66778 14504
rect 256786 14492 256792 14504
rect 256844 14492 256850 14544
rect 63218 14424 63224 14476
rect 63276 14464 63282 14476
rect 255498 14464 255504 14476
rect 63276 14436 255504 14464
rect 63276 14424 63282 14436
rect 255498 14424 255504 14436
rect 255556 14424 255562 14476
rect 102226 14356 102232 14408
rect 102284 14396 102290 14408
rect 269390 14396 269396 14408
rect 102284 14368 269396 14396
rect 102284 14356 102290 14368
rect 269390 14356 269396 14368
rect 269448 14356 269454 14408
rect 105722 14288 105728 14340
rect 105780 14328 105786 14340
rect 270586 14328 270592 14340
rect 105780 14300 270592 14328
rect 105780 14288 105786 14300
rect 270586 14288 270592 14300
rect 270644 14288 270650 14340
rect 109034 14220 109040 14272
rect 109092 14260 109098 14272
rect 272058 14260 272064 14272
rect 109092 14232 272064 14260
rect 109092 14220 109098 14232
rect 272058 14220 272064 14232
rect 272116 14220 272122 14272
rect 108114 13744 108120 13796
rect 108172 13784 108178 13796
rect 271966 13784 271972 13796
rect 108172 13756 271972 13784
rect 108172 13744 108178 13756
rect 271966 13744 271972 13756
rect 272024 13744 272030 13796
rect 404538 13744 404544 13796
rect 404596 13784 404602 13796
rect 497090 13784 497096 13796
rect 404596 13756 497096 13784
rect 404596 13744 404602 13756
rect 497090 13744 497096 13756
rect 497148 13744 497154 13796
rect 104066 13676 104072 13728
rect 104124 13716 104130 13728
rect 270678 13716 270684 13728
rect 104124 13688 270684 13716
rect 104124 13676 104130 13688
rect 270678 13676 270684 13688
rect 270736 13676 270742 13728
rect 405918 13676 405924 13728
rect 405976 13716 405982 13728
rect 500586 13716 500592 13728
rect 405976 13688 500592 13716
rect 405976 13676 405982 13688
rect 500586 13676 500592 13688
rect 500644 13676 500650 13728
rect 100754 13608 100760 13660
rect 100812 13648 100818 13660
rect 269298 13648 269304 13660
rect 100812 13620 269304 13648
rect 100812 13608 100818 13620
rect 269298 13608 269304 13620
rect 269356 13608 269362 13660
rect 407390 13608 407396 13660
rect 407448 13648 407454 13660
rect 503714 13648 503720 13660
rect 407448 13620 503720 13648
rect 407448 13608 407454 13620
rect 503714 13608 503720 13620
rect 503772 13608 503778 13660
rect 97442 13540 97448 13592
rect 97500 13580 97506 13592
rect 267918 13580 267924 13592
rect 97500 13552 267924 13580
rect 97500 13540 97506 13552
rect 267918 13540 267924 13552
rect 267976 13540 267982 13592
rect 408678 13540 408684 13592
rect 408736 13580 408742 13592
rect 507210 13580 507216 13592
rect 408736 13552 507216 13580
rect 408736 13540 408742 13552
rect 507210 13540 507216 13552
rect 507268 13540 507274 13592
rect 93946 13472 93952 13524
rect 94004 13512 94010 13524
rect 266538 13512 266544 13524
rect 94004 13484 266544 13512
rect 94004 13472 94010 13484
rect 266538 13472 266544 13484
rect 266596 13472 266602 13524
rect 410150 13472 410156 13524
rect 410208 13512 410214 13524
rect 511258 13512 511264 13524
rect 410208 13484 511264 13512
rect 410208 13472 410214 13484
rect 511258 13472 511264 13484
rect 511316 13472 511322 13524
rect 59354 13404 59360 13456
rect 59412 13444 59418 13456
rect 255406 13444 255412 13456
rect 59412 13416 255412 13444
rect 59412 13404 59418 13416
rect 255406 13404 255412 13416
rect 255464 13404 255470 13456
rect 411438 13404 411444 13456
rect 411496 13444 411502 13456
rect 514754 13444 514760 13456
rect 411496 13416 514760 13444
rect 411496 13404 411502 13416
rect 514754 13404 514760 13416
rect 514812 13404 514818 13456
rect 56042 13336 56048 13388
rect 56100 13376 56106 13388
rect 254026 13376 254032 13388
rect 56100 13348 254032 13376
rect 56100 13336 56106 13348
rect 254026 13336 254032 13348
rect 254084 13336 254090 13388
rect 414290 13336 414296 13388
rect 414348 13376 414354 13388
rect 521654 13376 521660 13388
rect 414348 13348 521660 13376
rect 414348 13336 414354 13348
rect 521654 13336 521660 13348
rect 521712 13336 521718 13388
rect 52546 13268 52552 13320
rect 52604 13308 52610 13320
rect 252738 13308 252744 13320
rect 52604 13280 252744 13308
rect 52604 13268 52610 13280
rect 252738 13268 252744 13280
rect 252796 13268 252802 13320
rect 414198 13268 414204 13320
rect 414256 13308 414262 13320
rect 525426 13308 525432 13320
rect 414256 13280 525432 13308
rect 414256 13268 414262 13280
rect 525426 13268 525432 13280
rect 525484 13268 525490 13320
rect 48498 13200 48504 13252
rect 48556 13240 48562 13252
rect 251266 13240 251272 13252
rect 48556 13212 251272 13240
rect 48556 13200 48562 13212
rect 251266 13200 251272 13212
rect 251324 13200 251330 13252
rect 417050 13200 417056 13252
rect 417108 13240 417114 13252
rect 532050 13240 532056 13252
rect 417108 13212 532056 13240
rect 417108 13200 417114 13212
rect 532050 13200 532056 13212
rect 532108 13200 532114 13252
rect 44266 13132 44272 13184
rect 44324 13172 44330 13184
rect 249978 13172 249984 13184
rect 44324 13144 249984 13172
rect 44324 13132 44330 13144
rect 249978 13132 249984 13144
rect 250036 13132 250042 13184
rect 422478 13132 422484 13184
rect 422536 13172 422542 13184
rect 546494 13172 546500 13184
rect 422536 13144 546500 13172
rect 422536 13132 422542 13144
rect 546494 13132 546500 13144
rect 546552 13132 546558 13184
rect 40218 13064 40224 13116
rect 40276 13104 40282 13116
rect 248506 13104 248512 13116
rect 40276 13076 248512 13104
rect 40276 13064 40282 13076
rect 248506 13064 248512 13076
rect 248564 13064 248570 13116
rect 429378 13064 429384 13116
rect 429436 13104 429442 13116
rect 567562 13104 567568 13116
rect 429436 13076 567568 13104
rect 429436 13064 429442 13076
rect 567562 13064 567568 13076
rect 567620 13064 567626 13116
rect 110414 12996 110420 13048
rect 110472 13036 110478 13048
rect 273346 13036 273352 13048
rect 110472 13008 273352 13036
rect 110472 12996 110478 13008
rect 273346 12996 273352 13008
rect 273404 12996 273410 13048
rect 403250 12996 403256 13048
rect 403308 13036 403314 13048
rect 493042 13036 493048 13048
rect 403308 13008 493048 13036
rect 403308 12996 403314 13008
rect 493042 12996 493048 13008
rect 493100 12996 493106 13048
rect 156138 12928 156144 12980
rect 156196 12968 156202 12980
rect 288618 12968 288624 12980
rect 156196 12940 288624 12968
rect 156196 12928 156202 12940
rect 288618 12928 288624 12940
rect 288676 12928 288682 12980
rect 390738 12928 390744 12980
rect 390796 12968 390802 12980
rect 454034 12968 454040 12980
rect 390796 12940 454040 12968
rect 390796 12928 390802 12940
rect 454034 12928 454040 12940
rect 454092 12928 454098 12980
rect 160094 12860 160100 12912
rect 160152 12900 160158 12912
rect 289998 12900 290004 12912
rect 160152 12872 290004 12900
rect 160152 12860 160158 12872
rect 289998 12860 290004 12872
rect 290056 12860 290062 12912
rect 219986 12384 219992 12436
rect 220044 12424 220050 12436
rect 310698 12424 310704 12436
rect 220044 12396 310704 12424
rect 220044 12384 220050 12396
rect 310698 12384 310704 12396
rect 310756 12384 310762 12436
rect 397638 12384 397644 12436
rect 397696 12424 397702 12436
rect 476482 12424 476488 12436
rect 397696 12396 476488 12424
rect 397696 12384 397702 12396
rect 476482 12384 476488 12396
rect 476540 12384 476546 12436
rect 216858 12316 216864 12368
rect 216916 12356 216922 12368
rect 309318 12356 309324 12368
rect 216916 12328 309324 12356
rect 216916 12316 216922 12328
rect 309318 12316 309324 12328
rect 309376 12316 309382 12368
rect 400490 12316 400496 12368
rect 400548 12356 400554 12368
rect 481726 12356 481732 12368
rect 400548 12328 481732 12356
rect 400548 12316 400554 12328
rect 481726 12316 481732 12328
rect 481784 12316 481790 12368
rect 213362 12248 213368 12300
rect 213420 12288 213426 12300
rect 308030 12288 308036 12300
rect 213420 12260 308036 12288
rect 213420 12248 213426 12260
rect 308030 12248 308036 12260
rect 308088 12248 308094 12300
rect 403158 12248 403164 12300
rect 403216 12288 403222 12300
rect 489914 12288 489920 12300
rect 403216 12260 489920 12288
rect 403216 12248 403222 12260
rect 489914 12248 489920 12260
rect 489972 12248 489978 12300
rect 209774 12180 209780 12232
rect 209832 12220 209838 12232
rect 306466 12220 306472 12232
rect 209832 12192 306472 12220
rect 209832 12180 209838 12192
rect 306466 12180 306472 12192
rect 306524 12180 306530 12232
rect 404446 12180 404452 12232
rect 404504 12220 404510 12232
rect 494698 12220 494704 12232
rect 404504 12192 494704 12220
rect 404504 12180 404510 12192
rect 494698 12180 494704 12192
rect 494756 12180 494762 12232
rect 206186 12112 206192 12164
rect 206244 12152 206250 12164
rect 305178 12152 305184 12164
rect 206244 12124 305184 12152
rect 206244 12112 206250 12124
rect 305178 12112 305184 12124
rect 305236 12112 305242 12164
rect 316218 12152 316224 12164
rect 316144 12124 316224 12152
rect 202690 12044 202696 12096
rect 202748 12084 202754 12096
rect 303798 12084 303804 12096
rect 202748 12056 303804 12084
rect 202748 12044 202754 12056
rect 303798 12044 303804 12056
rect 303856 12044 303862 12096
rect 145466 11976 145472 12028
rect 145524 12016 145530 12028
rect 284386 12016 284392 12028
rect 145524 11988 284392 12016
rect 145524 11976 145530 11988
rect 284386 11976 284392 11988
rect 284444 11976 284450 12028
rect 316144 11960 316172 12124
rect 316218 12112 316224 12124
rect 316276 12112 316282 12164
rect 418246 12112 418252 12164
rect 418304 12152 418310 12164
rect 534442 12152 534448 12164
rect 418304 12124 534448 12152
rect 418304 12112 418310 12124
rect 534442 12112 534448 12124
rect 534500 12112 534506 12164
rect 419718 12044 419724 12096
rect 419776 12084 419782 12096
rect 538214 12084 538220 12096
rect 419776 12056 538220 12084
rect 419776 12044 419782 12056
rect 538214 12044 538220 12056
rect 538272 12044 538278 12096
rect 421006 11976 421012 12028
rect 421064 12016 421070 12028
rect 541986 12016 541992 12028
rect 421064 11988 541992 12016
rect 421064 11976 421070 11988
rect 541986 11976 541992 11988
rect 542044 11976 542050 12028
rect 142154 11908 142160 11960
rect 142212 11948 142218 11960
rect 283006 11948 283012 11960
rect 142212 11920 283012 11948
rect 142212 11908 142218 11920
rect 283006 11908 283012 11920
rect 283064 11908 283070 11960
rect 316126 11908 316132 11960
rect 316184 11908 316190 11960
rect 421098 11908 421104 11960
rect 421156 11948 421162 11960
rect 545482 11948 545488 11960
rect 421156 11920 545488 11948
rect 421156 11908 421162 11920
rect 545482 11908 545488 11920
rect 545540 11908 545546 11960
rect 138842 11840 138848 11892
rect 138900 11880 138906 11892
rect 281718 11880 281724 11892
rect 138900 11852 281724 11880
rect 138900 11840 138906 11852
rect 281718 11840 281724 11852
rect 281776 11840 281782 11892
rect 422386 11840 422392 11892
rect 422444 11880 422450 11892
rect 547874 11880 547880 11892
rect 422444 11852 547880 11880
rect 422444 11840 422450 11852
rect 547874 11840 547880 11852
rect 547932 11840 547938 11892
rect 135254 11772 135260 11824
rect 135312 11812 135318 11824
rect 280338 11812 280344 11824
rect 135312 11784 280344 11812
rect 135312 11772 135318 11784
rect 280338 11772 280344 11784
rect 280396 11772 280402 11824
rect 423858 11772 423864 11824
rect 423916 11812 423922 11824
rect 551002 11812 551008 11824
rect 423916 11784 551008 11812
rect 423916 11772 423922 11784
rect 551002 11772 551008 11784
rect 551060 11772 551066 11824
rect 131298 11704 131304 11756
rect 131356 11744 131362 11756
rect 280430 11744 280436 11756
rect 131356 11716 280436 11744
rect 131356 11704 131362 11716
rect 280430 11704 280436 11716
rect 280488 11704 280494 11756
rect 425146 11704 425152 11756
rect 425204 11744 425210 11756
rect 554774 11744 554780 11756
rect 425204 11716 554780 11744
rect 425204 11704 425210 11716
rect 554774 11704 554780 11716
rect 554832 11704 554838 11756
rect 143534 11636 143540 11688
rect 143592 11676 143598 11688
rect 144730 11676 144736 11688
rect 143592 11648 144736 11676
rect 143592 11636 143598 11648
rect 144730 11636 144736 11648
rect 144788 11636 144794 11688
rect 223574 11636 223580 11688
rect 223632 11676 223638 11688
rect 310606 11676 310612 11688
rect 223632 11648 310612 11676
rect 223632 11636 223638 11648
rect 310606 11636 310612 11648
rect 310664 11636 310670 11688
rect 396442 11636 396448 11688
rect 396500 11676 396506 11688
rect 473446 11676 473452 11688
rect 396500 11648 473452 11676
rect 396500 11636 396506 11648
rect 473446 11636 473452 11648
rect 473504 11636 473510 11688
rect 226334 11568 226340 11620
rect 226392 11608 226398 11620
rect 312078 11608 312084 11620
rect 226392 11580 312084 11608
rect 226392 11568 226398 11580
rect 312078 11568 312084 11580
rect 312136 11568 312142 11620
rect 396350 11568 396356 11620
rect 396408 11608 396414 11620
rect 469858 11608 469864 11620
rect 396408 11580 469864 11608
rect 396408 11568 396414 11580
rect 469858 11568 469864 11580
rect 469916 11568 469922 11620
rect 231026 11500 231032 11552
rect 231084 11540 231090 11552
rect 313366 11540 313372 11552
rect 231084 11512 313372 11540
rect 231084 11500 231090 11512
rect 313366 11500 313372 11512
rect 313424 11500 313430 11552
rect 394786 11500 394792 11552
rect 394844 11540 394850 11552
rect 465626 11540 465632 11552
rect 394844 11512 465632 11540
rect 394844 11500 394850 11512
rect 465626 11500 465632 11512
rect 465684 11500 465690 11552
rect 173894 10956 173900 11008
rect 173952 10996 173958 11008
rect 294046 10996 294052 11008
rect 173952 10968 294052 10996
rect 173952 10956 173958 10968
rect 294046 10956 294052 10968
rect 294104 10956 294110 11008
rect 393406 10956 393412 11008
rect 393464 10996 393470 11008
rect 463970 10996 463976 11008
rect 393464 10968 463976 10996
rect 393464 10956 393470 10968
rect 463970 10956 463976 10968
rect 464028 10956 464034 11008
rect 170306 10888 170312 10940
rect 170364 10928 170370 10940
rect 292666 10928 292672 10940
rect 170364 10900 292672 10928
rect 170364 10888 170370 10900
rect 292666 10888 292672 10900
rect 292724 10888 292730 10940
rect 394694 10888 394700 10940
rect 394752 10928 394758 10940
rect 467466 10928 467472 10940
rect 394752 10900 467472 10928
rect 394752 10888 394758 10900
rect 467466 10888 467472 10900
rect 467524 10888 467530 10940
rect 167178 10820 167184 10872
rect 167236 10860 167242 10872
rect 291378 10860 291384 10872
rect 167236 10832 291384 10860
rect 167236 10820 167242 10832
rect 291378 10820 291384 10832
rect 291436 10820 291442 10872
rect 396258 10820 396264 10872
rect 396316 10860 396322 10872
rect 470594 10860 470600 10872
rect 396316 10832 470600 10860
rect 396316 10820 396322 10832
rect 470594 10820 470600 10832
rect 470652 10820 470658 10872
rect 163406 10752 163412 10804
rect 163464 10792 163470 10804
rect 289906 10792 289912 10804
rect 163464 10764 289912 10792
rect 163464 10752 163470 10764
rect 289906 10752 289912 10764
rect 289964 10752 289970 10804
rect 397546 10752 397552 10804
rect 397604 10792 397610 10804
rect 474090 10792 474096 10804
rect 397604 10764 474096 10792
rect 397604 10752 397610 10764
rect 474090 10752 474096 10764
rect 474148 10752 474154 10804
rect 158898 10684 158904 10736
rect 158956 10724 158962 10736
rect 288526 10724 288532 10736
rect 158956 10696 288532 10724
rect 158956 10684 158962 10696
rect 288526 10684 288532 10696
rect 288584 10684 288590 10736
rect 398926 10684 398932 10736
rect 398984 10724 398990 10736
rect 478138 10724 478144 10736
rect 398984 10696 478144 10724
rect 398984 10684 398990 10696
rect 478138 10684 478144 10696
rect 478196 10684 478202 10736
rect 155402 10616 155408 10668
rect 155460 10656 155466 10668
rect 287146 10656 287152 10668
rect 155460 10628 287152 10656
rect 155460 10616 155466 10628
rect 287146 10616 287152 10628
rect 287204 10616 287210 10668
rect 400398 10616 400404 10668
rect 400456 10656 400462 10668
rect 482370 10656 482376 10668
rect 400456 10628 482376 10656
rect 400456 10616 400462 10628
rect 482370 10616 482376 10628
rect 482428 10616 482434 10668
rect 89898 10548 89904 10600
rect 89956 10588 89962 10600
rect 265158 10588 265164 10600
rect 89956 10560 265164 10588
rect 89956 10548 89962 10560
rect 265158 10548 265164 10560
rect 265216 10548 265222 10600
rect 398834 10548 398840 10600
rect 398892 10588 398898 10600
rect 480530 10588 480536 10600
rect 398892 10560 480536 10588
rect 398892 10548 398898 10560
rect 480530 10548 480536 10560
rect 480588 10548 480594 10600
rect 86402 10480 86408 10532
rect 86460 10520 86466 10532
rect 263778 10520 263784 10532
rect 86460 10492 263784 10520
rect 86460 10480 86466 10492
rect 263778 10480 263784 10492
rect 263836 10480 263842 10532
rect 400306 10480 400312 10532
rect 400364 10520 400370 10532
rect 484026 10520 484032 10532
rect 400364 10492 484032 10520
rect 400364 10480 400370 10492
rect 484026 10480 484032 10492
rect 484084 10480 484090 10532
rect 83274 10412 83280 10464
rect 83332 10452 83338 10464
rect 262306 10452 262312 10464
rect 83332 10424 262312 10452
rect 83332 10412 83338 10424
rect 262306 10412 262312 10424
rect 262364 10412 262370 10464
rect 401686 10412 401692 10464
rect 401744 10452 401750 10464
rect 486418 10452 486424 10464
rect 401744 10424 486424 10452
rect 401744 10412 401750 10424
rect 486418 10412 486424 10424
rect 486476 10412 486482 10464
rect 79226 10344 79232 10396
rect 79284 10384 79290 10396
rect 262398 10384 262404 10396
rect 79284 10356 262404 10384
rect 79284 10344 79290 10356
rect 262398 10344 262404 10356
rect 262456 10344 262462 10396
rect 401778 10344 401784 10396
rect 401836 10384 401842 10396
rect 487154 10384 487160 10396
rect 401836 10356 487160 10384
rect 401836 10344 401842 10356
rect 487154 10344 487160 10356
rect 487212 10344 487218 10396
rect 75914 10276 75920 10328
rect 75972 10316 75978 10328
rect 261018 10316 261024 10328
rect 75972 10288 261024 10316
rect 75972 10276 75978 10288
rect 261018 10276 261024 10288
rect 261076 10276 261082 10328
rect 403066 10276 403072 10328
rect 403124 10316 403130 10328
rect 490650 10316 490656 10328
rect 403124 10288 490656 10316
rect 403124 10276 403130 10288
rect 490650 10276 490656 10288
rect 490708 10276 490714 10328
rect 176654 10208 176660 10260
rect 176712 10248 176718 10260
rect 295518 10248 295524 10260
rect 176712 10220 295524 10248
rect 176712 10208 176718 10220
rect 295518 10208 295524 10220
rect 295576 10208 295582 10260
rect 392118 10208 392124 10260
rect 392176 10248 392182 10260
rect 459922 10248 459928 10260
rect 392176 10220 459928 10248
rect 392176 10208 392182 10220
rect 459922 10208 459928 10220
rect 459980 10208 459986 10260
rect 180978 10140 180984 10192
rect 181036 10180 181042 10192
rect 297082 10180 297088 10192
rect 181036 10152 297088 10180
rect 181036 10140 181042 10152
rect 297082 10140 297088 10152
rect 297140 10140 297146 10192
rect 390646 10140 390652 10192
rect 390704 10180 390710 10192
rect 456886 10180 456892 10192
rect 390704 10152 456892 10180
rect 390704 10140 390710 10152
rect 456886 10140 456892 10152
rect 456944 10140 456950 10192
rect 184934 10072 184940 10124
rect 184992 10112 184998 10124
rect 298370 10112 298376 10124
rect 184992 10084 298376 10112
rect 184992 10072 184998 10084
rect 298370 10072 298376 10084
rect 298428 10072 298434 10124
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 222746 9596 222752 9648
rect 222804 9636 222810 9648
rect 310514 9636 310520 9648
rect 222804 9608 310520 9636
rect 222804 9596 222810 9608
rect 310514 9596 310520 9608
rect 310572 9596 310578 9648
rect 387886 9596 387892 9648
rect 387944 9636 387950 9648
rect 446214 9636 446220 9648
rect 387944 9608 446220 9636
rect 387944 9596 387950 9608
rect 446214 9596 446220 9608
rect 446272 9596 446278 9648
rect 219250 9528 219256 9580
rect 219308 9568 219314 9580
rect 309226 9568 309232 9580
rect 219308 9540 309232 9568
rect 219308 9528 219314 9540
rect 309226 9528 309232 9540
rect 309284 9528 309290 9580
rect 316034 9528 316040 9580
rect 316092 9568 316098 9580
rect 316310 9568 316316 9580
rect 316092 9540 316316 9568
rect 316092 9528 316098 9540
rect 316310 9528 316316 9540
rect 316368 9528 316374 9580
rect 389266 9528 389272 9580
rect 389324 9568 389330 9580
rect 449802 9568 449808 9580
rect 389324 9540 449808 9568
rect 389324 9528 389330 9540
rect 449802 9528 449808 9540
rect 449860 9528 449866 9580
rect 215662 9460 215668 9512
rect 215720 9500 215726 9512
rect 307938 9500 307944 9512
rect 215720 9472 307944 9500
rect 215720 9460 215726 9472
rect 307938 9460 307944 9472
rect 307996 9460 308002 9512
rect 315942 9460 315948 9512
rect 316000 9500 316006 9512
rect 316218 9500 316224 9512
rect 316000 9472 316224 9500
rect 316000 9460 316006 9472
rect 316218 9460 316224 9472
rect 316276 9460 316282 9512
rect 389358 9460 389364 9512
rect 389416 9500 389422 9512
rect 453298 9500 453304 9512
rect 389416 9472 453304 9500
rect 389416 9460 389422 9472
rect 453298 9460 453304 9472
rect 453356 9460 453362 9512
rect 137646 9392 137652 9444
rect 137704 9432 137710 9444
rect 281626 9432 281632 9444
rect 137704 9404 281632 9432
rect 137704 9392 137710 9404
rect 281626 9392 281632 9404
rect 281684 9392 281690 9444
rect 422294 9392 422300 9444
rect 422352 9432 422358 9444
rect 549070 9432 549076 9444
rect 422352 9404 549076 9432
rect 422352 9392 422358 9404
rect 549070 9392 549076 9404
rect 549128 9392 549134 9444
rect 37182 9324 37188 9376
rect 37240 9364 37246 9376
rect 247126 9364 247132 9376
rect 37240 9336 247132 9364
rect 37240 9324 37246 9336
rect 247126 9324 247132 9336
rect 247184 9324 247190 9376
rect 277118 9324 277124 9376
rect 277176 9364 277182 9376
rect 330018 9364 330024 9376
rect 277176 9336 330024 9364
rect 277176 9324 277182 9336
rect 330018 9324 330024 9336
rect 330076 9324 330082 9376
rect 423766 9324 423772 9376
rect 423824 9364 423830 9376
rect 552658 9364 552664 9376
rect 423824 9336 552664 9364
rect 423824 9324 423830 9336
rect 552658 9324 552664 9336
rect 552716 9324 552722 9376
rect 33594 9256 33600 9308
rect 33652 9296 33658 9308
rect 245930 9296 245936 9308
rect 33652 9268 245936 9296
rect 33652 9256 33658 9268
rect 245930 9256 245936 9268
rect 245988 9256 245994 9308
rect 262950 9256 262956 9308
rect 263008 9296 263014 9308
rect 324590 9296 324596 9308
rect 263008 9268 324596 9296
rect 263008 9256 263014 9268
rect 324590 9256 324596 9268
rect 324648 9256 324654 9308
rect 425054 9256 425060 9308
rect 425112 9296 425118 9308
rect 556154 9296 556160 9308
rect 425112 9268 556160 9296
rect 425112 9256 425118 9268
rect 556154 9256 556160 9268
rect 556212 9256 556218 9308
rect 30098 9188 30104 9240
rect 30156 9228 30162 9240
rect 244366 9228 244372 9240
rect 30156 9200 244372 9228
rect 30156 9188 30162 9200
rect 244366 9188 244372 9200
rect 244424 9188 244430 9240
rect 259454 9188 259460 9240
rect 259512 9228 259518 9240
rect 323118 9228 323124 9240
rect 259512 9200 323124 9228
rect 259512 9188 259518 9200
rect 323118 9188 323124 9200
rect 323176 9188 323182 9240
rect 426526 9188 426532 9240
rect 426584 9228 426590 9240
rect 559742 9228 559748 9240
rect 426584 9200 559748 9228
rect 426584 9188 426590 9200
rect 559742 9188 559748 9200
rect 559800 9188 559806 9240
rect 26510 9120 26516 9172
rect 26568 9160 26574 9172
rect 242986 9160 242992 9172
rect 26568 9132 242992 9160
rect 26568 9120 26574 9132
rect 242986 9120 242992 9132
rect 243044 9120 243050 9172
rect 255866 9120 255872 9172
rect 255924 9160 255930 9172
rect 321830 9160 321836 9172
rect 255924 9132 321836 9160
rect 255924 9120 255930 9132
rect 321830 9120 321836 9132
rect 321888 9120 321894 9172
rect 427998 9120 428004 9172
rect 428056 9160 428062 9172
rect 563238 9160 563244 9172
rect 428056 9132 563244 9160
rect 428056 9120 428062 9132
rect 563238 9120 563244 9132
rect 563296 9120 563302 9172
rect 21818 9052 21824 9104
rect 21876 9092 21882 9104
rect 241698 9092 241704 9104
rect 21876 9064 241704 9092
rect 21876 9052 21882 9064
rect 241698 9052 241704 9064
rect 241756 9052 241762 9104
rect 252370 9052 252376 9104
rect 252428 9092 252434 9104
rect 321738 9092 321744 9104
rect 252428 9064 321744 9092
rect 252428 9052 252434 9064
rect 321738 9052 321744 9064
rect 321796 9052 321802 9104
rect 429286 9052 429292 9104
rect 429344 9092 429350 9104
rect 566826 9092 566832 9104
rect 429344 9064 566832 9092
rect 429344 9052 429350 9064
rect 566826 9052 566832 9064
rect 566884 9052 566890 9104
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 237466 9024 237472 9036
rect 8812 8996 237472 9024
rect 8812 8984 8818 8996
rect 237466 8984 237472 8996
rect 237524 8984 237530 9036
rect 242066 8984 242072 9036
rect 242124 9024 242130 9036
rect 317690 9024 317696 9036
rect 242124 8996 317696 9024
rect 242124 8984 242130 8996
rect 317690 8984 317696 8996
rect 317748 8984 317754 9036
rect 430758 8984 430764 9036
rect 430816 9024 430822 9036
rect 570322 9024 570328 9036
rect 430816 8996 570328 9024
rect 430816 8984 430822 8996
rect 570322 8984 570328 8996
rect 570380 8984 570386 9036
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 236086 8956 236092 8968
rect 4120 8928 236092 8956
rect 4120 8916 4126 8928
rect 236086 8916 236092 8928
rect 236144 8916 236150 8968
rect 238110 8916 238116 8968
rect 238168 8956 238174 8968
rect 316402 8956 316408 8968
rect 238168 8928 316408 8956
rect 238168 8916 238174 8928
rect 316402 8916 316408 8928
rect 316460 8916 316466 8968
rect 430666 8916 430672 8968
rect 430724 8956 430730 8968
rect 573910 8956 573916 8968
rect 430724 8928 573916 8956
rect 430724 8916 430730 8928
rect 573910 8916 573916 8928
rect 573968 8916 573974 8968
rect 226426 8848 226432 8900
rect 226484 8888 226490 8900
rect 311986 8888 311992 8900
rect 226484 8860 311992 8888
rect 226484 8848 226490 8860
rect 311986 8848 311992 8860
rect 312044 8848 312050 8900
rect 386690 8848 386696 8900
rect 386748 8888 386754 8900
rect 442626 8888 442632 8900
rect 386748 8860 442632 8888
rect 386748 8848 386754 8860
rect 442626 8848 442632 8860
rect 442684 8848 442690 8900
rect 229830 8780 229836 8832
rect 229888 8820 229894 8832
rect 313274 8820 313280 8832
rect 229888 8792 313280 8820
rect 229888 8780 229894 8792
rect 313274 8780 313280 8792
rect 313332 8780 313338 8832
rect 385126 8780 385132 8832
rect 385184 8820 385190 8832
rect 439130 8820 439136 8832
rect 385184 8792 439136 8820
rect 385184 8780 385190 8792
rect 439130 8780 439136 8792
rect 439188 8780 439194 8832
rect 233418 8712 233424 8764
rect 233476 8752 233482 8764
rect 314838 8752 314844 8764
rect 233476 8724 314844 8752
rect 233476 8712 233482 8724
rect 314838 8712 314844 8724
rect 314896 8712 314902 8764
rect 383838 8712 383844 8764
rect 383896 8752 383902 8764
rect 435542 8752 435548 8764
rect 383896 8724 435548 8752
rect 383896 8712 383902 8724
rect 435542 8712 435548 8724
rect 435600 8712 435606 8764
rect 183738 8236 183744 8288
rect 183796 8276 183802 8288
rect 296898 8276 296904 8288
rect 183796 8248 296904 8276
rect 183796 8236 183802 8248
rect 296898 8236 296904 8248
rect 296956 8236 296962 8288
rect 404354 8236 404360 8288
rect 404412 8276 404418 8288
rect 495894 8276 495900 8288
rect 404412 8248 495900 8276
rect 404412 8236 404418 8248
rect 495894 8236 495900 8248
rect 495952 8236 495958 8288
rect 180242 8168 180248 8220
rect 180300 8208 180306 8220
rect 296990 8208 296996 8220
rect 180300 8180 296996 8208
rect 180300 8168 180306 8180
rect 296990 8168 296996 8180
rect 297048 8168 297054 8220
rect 405826 8168 405832 8220
rect 405884 8208 405890 8220
rect 499390 8208 499396 8220
rect 405884 8180 499396 8208
rect 405884 8168 405890 8180
rect 499390 8168 499396 8180
rect 499448 8168 499454 8220
rect 176746 8100 176752 8152
rect 176804 8140 176810 8152
rect 295426 8140 295432 8152
rect 176804 8112 295432 8140
rect 176804 8100 176810 8112
rect 295426 8100 295432 8112
rect 295484 8100 295490 8152
rect 407298 8100 407304 8152
rect 407356 8140 407362 8152
rect 502978 8140 502984 8152
rect 407356 8112 502984 8140
rect 407356 8100 407362 8112
rect 502978 8100 502984 8112
rect 503036 8100 503042 8152
rect 173066 8032 173072 8084
rect 173124 8072 173130 8084
rect 294230 8072 294236 8084
rect 173124 8044 294236 8072
rect 173124 8032 173130 8044
rect 294230 8032 294236 8044
rect 294288 8032 294294 8084
rect 408586 8032 408592 8084
rect 408644 8072 408650 8084
rect 506474 8072 506480 8084
rect 408644 8044 506480 8072
rect 408644 8032 408650 8044
rect 506474 8032 506480 8044
rect 506532 8032 506538 8084
rect 169570 7964 169576 8016
rect 169628 8004 169634 8016
rect 292574 8004 292580 8016
rect 169628 7976 292580 8004
rect 169628 7964 169634 7976
rect 292574 7964 292580 7976
rect 292632 7964 292638 8016
rect 409966 7964 409972 8016
rect 410024 8004 410030 8016
rect 510062 8004 510068 8016
rect 410024 7976 510068 8004
rect 410024 7964 410030 7976
rect 510062 7964 510068 7976
rect 510120 7964 510126 8016
rect 162486 7896 162492 7948
rect 162544 7936 162550 7948
rect 289814 7936 289820 7948
rect 162544 7908 289820 7936
rect 162544 7896 162550 7908
rect 289814 7896 289820 7908
rect 289872 7896 289878 7948
rect 290734 7896 290740 7948
rect 290792 7936 290798 7948
rect 320358 7936 320364 7948
rect 290792 7908 320364 7936
rect 290792 7896 290798 7908
rect 320358 7896 320364 7908
rect 320416 7896 320422 7948
rect 410058 7896 410064 7948
rect 410116 7936 410122 7948
rect 513558 7936 513564 7948
rect 410116 7908 513564 7936
rect 410116 7896 410122 7908
rect 513558 7896 513564 7908
rect 513616 7896 513622 7948
rect 157794 7828 157800 7880
rect 157852 7868 157858 7880
rect 288434 7868 288440 7880
rect 157852 7840 288440 7868
rect 157852 7828 157858 7840
rect 288434 7828 288440 7840
rect 288492 7828 288498 7880
rect 288526 7828 288532 7880
rect 288584 7868 288590 7880
rect 328546 7868 328552 7880
rect 288584 7840 328552 7868
rect 288584 7828 288590 7840
rect 328546 7828 328552 7840
rect 328604 7828 328610 7880
rect 411346 7828 411352 7880
rect 411404 7868 411410 7880
rect 517146 7868 517152 7880
rect 411404 7840 517152 7868
rect 411404 7828 411410 7840
rect 517146 7828 517152 7840
rect 517204 7828 517210 7880
rect 130562 7760 130568 7812
rect 130620 7800 130626 7812
rect 278958 7800 278964 7812
rect 130620 7772 278964 7800
rect 130620 7760 130626 7772
rect 278958 7760 278964 7772
rect 279016 7760 279022 7812
rect 286594 7760 286600 7812
rect 286652 7800 286658 7812
rect 332686 7800 332692 7812
rect 286652 7772 332692 7800
rect 286652 7760 286658 7772
rect 332686 7760 332692 7772
rect 332744 7760 332750 7812
rect 412726 7760 412732 7812
rect 412784 7800 412790 7812
rect 520734 7800 520740 7812
rect 412784 7772 520740 7800
rect 412784 7760 412790 7772
rect 520734 7760 520740 7772
rect 520792 7760 520798 7812
rect 126974 7692 126980 7744
rect 127032 7732 127038 7744
rect 277578 7732 277584 7744
rect 127032 7704 277584 7732
rect 127032 7692 127038 7704
rect 277578 7692 277584 7704
rect 277636 7692 277642 7744
rect 283098 7692 283104 7744
rect 283156 7732 283162 7744
rect 331490 7732 331496 7744
rect 283156 7704 331496 7732
rect 283156 7692 283162 7704
rect 331490 7692 331496 7704
rect 331548 7692 331554 7744
rect 414106 7692 414112 7744
rect 414164 7732 414170 7744
rect 524230 7732 524236 7744
rect 414164 7704 524236 7732
rect 414164 7692 414170 7704
rect 524230 7692 524236 7704
rect 524288 7692 524294 7744
rect 128170 7624 128176 7676
rect 128228 7664 128234 7676
rect 278866 7664 278872 7676
rect 128228 7636 278872 7664
rect 128228 7624 128234 7636
rect 278866 7624 278872 7636
rect 278924 7624 278930 7676
rect 279510 7624 279516 7676
rect 279568 7664 279574 7676
rect 329926 7664 329932 7676
rect 279568 7636 329932 7664
rect 279568 7624 279574 7636
rect 329926 7624 329932 7636
rect 329984 7624 329990 7676
rect 415486 7624 415492 7676
rect 415544 7664 415550 7676
rect 527818 7664 527824 7676
rect 415544 7636 527824 7664
rect 415544 7624 415550 7636
rect 527818 7624 527824 7636
rect 527876 7624 527882 7676
rect 69106 7556 69112 7608
rect 69164 7596 69170 7608
rect 258074 7596 258080 7608
rect 69164 7568 258080 7596
rect 69164 7556 69170 7568
rect 258074 7556 258080 7568
rect 258132 7556 258138 7608
rect 272426 7556 272432 7608
rect 272484 7596 272490 7608
rect 328638 7596 328644 7608
rect 272484 7568 328644 7596
rect 272484 7556 272490 7568
rect 328638 7556 328644 7568
rect 328696 7556 328702 7608
rect 416958 7556 416964 7608
rect 417016 7596 417022 7608
rect 531314 7596 531320 7608
rect 417016 7568 531320 7596
rect 417016 7556 417022 7568
rect 531314 7556 531320 7568
rect 531372 7556 531378 7608
rect 187326 7488 187332 7540
rect 187384 7528 187390 7540
rect 298278 7528 298284 7540
rect 187384 7500 298284 7528
rect 187384 7488 187390 7500
rect 298278 7488 298284 7500
rect 298336 7488 298342 7540
rect 402974 7488 402980 7540
rect 403032 7528 403038 7540
rect 492306 7528 492312 7540
rect 403032 7500 492312 7528
rect 403032 7488 403038 7500
rect 492306 7488 492312 7500
rect 492364 7488 492370 7540
rect 190822 7420 190828 7472
rect 190880 7460 190886 7472
rect 299566 7460 299572 7472
rect 190880 7432 299572 7460
rect 190880 7420 190886 7432
rect 299566 7420 299572 7432
rect 299624 7420 299630 7472
rect 401594 7420 401600 7472
rect 401652 7460 401658 7472
rect 488810 7460 488816 7472
rect 401652 7432 488816 7460
rect 401652 7420 401658 7432
rect 488810 7420 488816 7432
rect 488868 7420 488874 7472
rect 194410 7352 194416 7404
rect 194468 7392 194474 7404
rect 300946 7392 300952 7404
rect 194468 7364 300952 7392
rect 194468 7352 194474 7364
rect 300946 7352 300952 7364
rect 301004 7352 301010 7404
rect 400214 7352 400220 7404
rect 400272 7392 400278 7404
rect 485222 7392 485228 7404
rect 400272 7364 485228 7392
rect 400272 7352 400278 7364
rect 485222 7352 485228 7364
rect 485280 7352 485286 7404
rect 62022 6808 62028 6860
rect 62080 6848 62086 6860
rect 255314 6848 255320 6860
rect 62080 6820 255320 6848
rect 62080 6808 62086 6820
rect 255314 6808 255320 6820
rect 255372 6808 255378 6860
rect 271230 6808 271236 6860
rect 271288 6848 271294 6860
rect 327166 6848 327172 6860
rect 271288 6820 327172 6848
rect 271288 6808 271294 6820
rect 327166 6808 327172 6820
rect 327224 6808 327230 6860
rect 387794 6808 387800 6860
rect 387852 6848 387858 6860
rect 448606 6848 448612 6860
rect 387852 6820 448612 6848
rect 387852 6808 387858 6820
rect 448606 6808 448612 6820
rect 448664 6808 448670 6860
rect 58434 6740 58440 6792
rect 58492 6780 58498 6792
rect 253934 6780 253940 6792
rect 58492 6752 253940 6780
rect 58492 6740 58498 6752
rect 253934 6740 253940 6752
rect 253992 6740 253998 6792
rect 268838 6740 268844 6792
rect 268896 6780 268902 6792
rect 327258 6780 327264 6792
rect 268896 6752 327264 6780
rect 268896 6740 268902 6752
rect 327258 6740 327264 6752
rect 327316 6740 327322 6792
rect 389174 6740 389180 6792
rect 389232 6780 389238 6792
rect 452102 6780 452108 6792
rect 389232 6752 452108 6780
rect 389232 6740 389238 6752
rect 452102 6740 452108 6752
rect 452160 6740 452166 6792
rect 54938 6672 54944 6724
rect 54996 6712 55002 6724
rect 252554 6712 252560 6724
rect 54996 6684 252560 6712
rect 54996 6672 55002 6684
rect 252554 6672 252560 6684
rect 252612 6672 252618 6724
rect 265342 6672 265348 6724
rect 265400 6712 265406 6724
rect 325878 6712 325884 6724
rect 265400 6684 325884 6712
rect 265400 6672 265406 6684
rect 325878 6672 325884 6684
rect 325936 6672 325942 6724
rect 390554 6672 390560 6724
rect 390612 6712 390618 6724
rect 455690 6712 455696 6724
rect 390612 6684 455696 6712
rect 390612 6672 390618 6684
rect 455690 6672 455696 6684
rect 455748 6672 455754 6724
rect 51350 6604 51356 6656
rect 51408 6644 51414 6656
rect 252646 6644 252652 6656
rect 51408 6616 252652 6644
rect 51408 6604 51414 6616
rect 252646 6604 252652 6616
rect 252704 6604 252710 6656
rect 261754 6604 261760 6656
rect 261812 6644 261818 6656
rect 324498 6644 324504 6656
rect 261812 6616 324504 6644
rect 261812 6604 261818 6616
rect 324498 6604 324504 6616
rect 324556 6604 324562 6656
rect 392026 6604 392032 6656
rect 392084 6644 392090 6656
rect 459186 6644 459192 6656
rect 392084 6616 459192 6644
rect 392084 6604 392090 6616
rect 459186 6604 459192 6616
rect 459244 6604 459250 6656
rect 47854 6536 47860 6588
rect 47912 6576 47918 6588
rect 251174 6576 251180 6588
rect 47912 6548 251180 6576
rect 47912 6536 47918 6548
rect 251174 6536 251180 6548
rect 251232 6536 251238 6588
rect 258258 6536 258264 6588
rect 258316 6576 258322 6588
rect 323026 6576 323032 6588
rect 258316 6548 323032 6576
rect 258316 6536 258322 6548
rect 323026 6536 323032 6548
rect 323084 6536 323090 6588
rect 393314 6536 393320 6588
rect 393372 6576 393378 6588
rect 462774 6576 462780 6588
rect 393372 6548 462780 6576
rect 393372 6536 393378 6548
rect 462774 6536 462780 6548
rect 462832 6536 462838 6588
rect 17034 6468 17040 6520
rect 17092 6508 17098 6520
rect 240318 6508 240324 6520
rect 17092 6480 240324 6508
rect 17092 6468 17098 6480
rect 240318 6468 240324 6480
rect 240376 6468 240382 6520
rect 254670 6468 254676 6520
rect 254728 6508 254734 6520
rect 321646 6508 321652 6520
rect 254728 6480 321652 6508
rect 254728 6468 254734 6480
rect 321646 6468 321652 6480
rect 321704 6468 321710 6520
rect 383746 6468 383752 6520
rect 383804 6508 383810 6520
rect 433978 6508 433984 6520
rect 383804 6480 412634 6508
rect 383804 6468 383810 6480
rect 12342 6400 12348 6452
rect 12400 6440 12406 6452
rect 238938 6440 238944 6452
rect 12400 6412 238944 6440
rect 12400 6400 12406 6412
rect 238938 6400 238944 6412
rect 238996 6400 239002 6452
rect 251174 6400 251180 6452
rect 251232 6440 251238 6452
rect 320266 6440 320272 6452
rect 251232 6412 320272 6440
rect 251232 6400 251238 6412
rect 320266 6400 320272 6412
rect 320324 6400 320330 6452
rect 412606 6440 412634 6480
rect 431926 6480 433984 6508
rect 431926 6440 431954 6480
rect 433978 6468 433984 6480
rect 434036 6468 434042 6520
rect 434070 6468 434076 6520
rect 434128 6508 434134 6520
rect 518342 6508 518348 6520
rect 434128 6480 518348 6508
rect 434128 6468 434134 6480
rect 518342 6468 518348 6480
rect 518400 6468 518406 6520
rect 562042 6440 562048 6452
rect 412606 6412 431954 6440
rect 433352 6412 562048 6440
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 237374 6372 237380 6384
rect 7708 6344 237380 6372
rect 7708 6332 7714 6344
rect 237374 6332 237380 6344
rect 237432 6332 237438 6384
rect 239306 6332 239312 6384
rect 239364 6372 239370 6384
rect 316126 6372 316132 6384
rect 239364 6344 316132 6372
rect 239364 6332 239370 6344
rect 316126 6332 316132 6344
rect 316184 6332 316190 6384
rect 379698 6332 379704 6384
rect 379756 6372 379762 6384
rect 424962 6372 424968 6384
rect 379756 6344 424968 6372
rect 379756 6332 379762 6344
rect 424962 6332 424968 6344
rect 425020 6332 425026 6384
rect 427906 6332 427912 6384
rect 427964 6372 427970 6384
rect 433352 6372 433380 6412
rect 562042 6400 562048 6412
rect 562100 6400 562106 6452
rect 427964 6344 433380 6372
rect 427964 6332 427970 6344
rect 436738 6332 436744 6384
rect 436796 6372 436802 6384
rect 565630 6372 565636 6384
rect 436796 6344 565636 6372
rect 436796 6332 436802 6344
rect 565630 6332 565636 6344
rect 565688 6332 565694 6384
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 234706 6304 234712 6316
rect 2924 6276 234712 6304
rect 2924 6264 2930 6276
rect 234706 6264 234712 6276
rect 234764 6264 234770 6316
rect 240502 6264 240508 6316
rect 240560 6304 240566 6316
rect 317598 6304 317604 6316
rect 240560 6276 317604 6304
rect 240560 6264 240566 6276
rect 317598 6264 317604 6276
rect 317656 6264 317662 6316
rect 380986 6264 380992 6316
rect 381044 6304 381050 6316
rect 427262 6304 427268 6316
rect 381044 6276 427268 6304
rect 381044 6264 381050 6276
rect 427262 6264 427268 6276
rect 427320 6264 427326 6316
rect 429194 6264 429200 6316
rect 429252 6304 429258 6316
rect 569126 6304 569132 6316
rect 429252 6276 569132 6304
rect 429252 6264 429258 6276
rect 569126 6264 569132 6276
rect 569184 6264 569190 6316
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 234798 6236 234804 6248
rect 1728 6208 234804 6236
rect 1728 6196 1734 6208
rect 234798 6196 234804 6208
rect 234856 6196 234862 6248
rect 235810 6196 235816 6248
rect 235868 6236 235874 6248
rect 314746 6236 314752 6248
rect 235868 6208 314752 6236
rect 235868 6196 235874 6208
rect 314746 6196 314752 6208
rect 314804 6196 314810 6248
rect 381078 6196 381084 6248
rect 381136 6236 381142 6248
rect 428458 6236 428464 6248
rect 381136 6208 428464 6236
rect 381136 6196 381142 6208
rect 428458 6196 428464 6208
rect 428516 6196 428522 6248
rect 430574 6196 430580 6248
rect 430632 6236 430638 6248
rect 572714 6236 572720 6248
rect 430632 6208 572720 6236
rect 430632 6196 430638 6208
rect 572714 6196 572720 6208
rect 572772 6196 572778 6248
rect 566 6128 572 6180
rect 624 6168 630 6180
rect 234614 6168 234620 6180
rect 624 6140 234620 6168
rect 624 6128 630 6140
rect 234614 6128 234620 6140
rect 234672 6128 234678 6180
rect 237006 6128 237012 6180
rect 237064 6168 237070 6180
rect 316034 6168 316040 6180
rect 237064 6140 316040 6168
rect 237064 6128 237070 6140
rect 316034 6128 316040 6140
rect 316092 6128 316098 6180
rect 432046 6128 432052 6180
rect 432104 6168 432110 6180
rect 576302 6168 576308 6180
rect 432104 6140 576308 6168
rect 432104 6128 432110 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 65518 6060 65524 6112
rect 65576 6100 65582 6112
rect 256694 6100 256700 6112
rect 65576 6072 256700 6100
rect 65576 6060 65582 6072
rect 256694 6060 256700 6072
rect 256752 6060 256758 6112
rect 285398 6060 285404 6112
rect 285456 6100 285462 6112
rect 332778 6100 332784 6112
rect 285456 6072 332784 6100
rect 285456 6060 285462 6072
rect 332778 6060 332784 6072
rect 332836 6060 332842 6112
rect 386506 6060 386512 6112
rect 386564 6100 386570 6112
rect 445018 6100 445024 6112
rect 386564 6072 445024 6100
rect 386564 6060 386570 6072
rect 445018 6060 445024 6072
rect 445076 6060 445082 6112
rect 136450 5992 136456 6044
rect 136508 6032 136514 6044
rect 281534 6032 281540 6044
rect 136508 6004 281540 6032
rect 136508 5992 136514 6004
rect 281534 5992 281540 6004
rect 281592 5992 281598 6044
rect 288986 5992 288992 6044
rect 289044 6032 289050 6044
rect 334066 6032 334072 6044
rect 289044 6004 334072 6032
rect 289044 5992 289050 6004
rect 334066 5992 334072 6004
rect 334124 5992 334130 6044
rect 386598 5992 386604 6044
rect 386656 6032 386662 6044
rect 441522 6032 441528 6044
rect 386656 6004 441528 6032
rect 386656 5992 386662 6004
rect 441522 5992 441528 6004
rect 441580 5992 441586 6044
rect 140038 5924 140044 5976
rect 140096 5964 140102 5976
rect 282914 5964 282920 5976
rect 140096 5936 282920 5964
rect 140096 5924 140102 5936
rect 282914 5924 282920 5936
rect 282972 5924 282978 5976
rect 309870 5924 309876 5976
rect 309928 5964 309934 5976
rect 334158 5964 334164 5976
rect 309928 5936 334164 5964
rect 309928 5924 309934 5936
rect 334158 5924 334164 5936
rect 334216 5924 334222 5976
rect 385034 5924 385040 5976
rect 385092 5964 385098 5976
rect 437934 5964 437940 5976
rect 385092 5936 437940 5964
rect 385092 5924 385098 5936
rect 437934 5924 437940 5936
rect 437992 5924 437998 5976
rect 234614 5856 234620 5908
rect 234672 5896 234678 5908
rect 262858 5896 262864 5908
rect 234672 5868 262864 5896
rect 234672 5856 234678 5868
rect 262858 5856 262864 5868
rect 262916 5856 262922 5908
rect 382550 5856 382556 5908
rect 382608 5896 382614 5908
rect 430850 5896 430856 5908
rect 382608 5868 430856 5896
rect 382608 5856 382614 5868
rect 430850 5856 430856 5868
rect 430908 5856 430914 5908
rect 382458 5788 382464 5840
rect 382516 5828 382522 5840
rect 432046 5828 432052 5840
rect 382516 5800 432052 5828
rect 382516 5788 382522 5800
rect 432046 5788 432052 5800
rect 432104 5788 432110 5840
rect 427814 5720 427820 5772
rect 427872 5760 427878 5772
rect 436738 5760 436744 5772
rect 427872 5732 436744 5760
rect 427872 5720 427878 5732
rect 436738 5720 436744 5732
rect 436796 5720 436802 5772
rect 210970 5448 210976 5500
rect 211028 5488 211034 5500
rect 306374 5488 306380 5500
rect 211028 5460 306380 5488
rect 211028 5448 211034 5460
rect 306374 5448 306380 5460
rect 306432 5448 306438 5500
rect 407206 5448 407212 5500
rect 407264 5488 407270 5500
rect 505370 5488 505376 5500
rect 407264 5460 505376 5488
rect 407264 5448 407270 5460
rect 505370 5448 505376 5460
rect 505428 5448 505434 5500
rect 85666 5380 85672 5432
rect 85724 5420 85730 5432
rect 149698 5420 149704 5432
rect 85724 5392 149704 5420
rect 85724 5380 85730 5392
rect 149698 5380 149704 5392
rect 149756 5380 149762 5432
rect 207382 5380 207388 5432
rect 207440 5420 207446 5432
rect 305086 5420 305092 5432
rect 207440 5392 305092 5420
rect 207440 5380 207446 5392
rect 305086 5380 305092 5392
rect 305144 5380 305150 5432
rect 324406 5380 324412 5432
rect 324464 5420 324470 5432
rect 345290 5420 345296 5432
rect 324464 5392 345296 5420
rect 324464 5380 324470 5392
rect 345290 5380 345296 5392
rect 345348 5380 345354 5432
rect 408494 5380 408500 5432
rect 408552 5420 408558 5432
rect 508866 5420 508872 5432
rect 408552 5392 508872 5420
rect 408552 5380 408558 5392
rect 508866 5380 508872 5392
rect 508924 5380 508930 5432
rect 89162 5312 89168 5364
rect 89220 5352 89226 5364
rect 153838 5352 153844 5364
rect 89220 5324 153844 5352
rect 89220 5312 89226 5324
rect 153838 5312 153844 5324
rect 153896 5312 153902 5364
rect 203886 5312 203892 5364
rect 203944 5352 203950 5364
rect 303614 5352 303620 5364
rect 203944 5324 303620 5352
rect 203944 5312 203950 5324
rect 303614 5312 303620 5324
rect 303672 5312 303678 5364
rect 317322 5312 317328 5364
rect 317380 5352 317386 5364
rect 343726 5352 343732 5364
rect 317380 5324 343732 5352
rect 317380 5312 317386 5324
rect 343726 5312 343732 5324
rect 343784 5312 343790 5364
rect 409874 5312 409880 5364
rect 409932 5352 409938 5364
rect 512454 5352 512460 5364
rect 409932 5324 512460 5352
rect 409932 5312 409938 5324
rect 512454 5312 512460 5324
rect 512512 5312 512518 5364
rect 78582 5244 78588 5296
rect 78640 5284 78646 5296
rect 145558 5284 145564 5296
rect 78640 5256 145564 5284
rect 78640 5244 78646 5256
rect 145558 5244 145564 5256
rect 145616 5244 145622 5296
rect 196802 5244 196808 5296
rect 196860 5284 196866 5296
rect 302234 5284 302240 5296
rect 196860 5256 302240 5284
rect 196860 5244 196866 5256
rect 302234 5244 302240 5256
rect 302292 5244 302298 5296
rect 313826 5244 313832 5296
rect 313884 5284 313890 5296
rect 342346 5284 342352 5296
rect 313884 5256 342352 5284
rect 313884 5244 313890 5256
rect 342346 5244 342352 5256
rect 342404 5244 342410 5296
rect 411254 5244 411260 5296
rect 411312 5284 411318 5296
rect 515950 5284 515956 5296
rect 411312 5256 515956 5284
rect 411312 5244 411318 5256
rect 515950 5244 515956 5256
rect 516008 5244 516014 5296
rect 96246 5176 96252 5228
rect 96304 5216 96310 5228
rect 163498 5216 163504 5228
rect 96304 5188 163504 5216
rect 96304 5176 96310 5188
rect 163498 5176 163504 5188
rect 163556 5176 163562 5228
rect 193214 5176 193220 5228
rect 193272 5216 193278 5228
rect 300854 5216 300860 5228
rect 193272 5188 300860 5216
rect 193272 5176 193278 5188
rect 300854 5176 300860 5188
rect 300912 5176 300918 5228
rect 310238 5176 310244 5228
rect 310296 5216 310302 5228
rect 341058 5216 341064 5228
rect 310296 5188 341064 5216
rect 310296 5176 310302 5188
rect 341058 5176 341064 5188
rect 341116 5176 341122 5228
rect 367278 5176 367284 5228
rect 367336 5216 367342 5228
rect 387150 5216 387156 5228
rect 367336 5188 387156 5216
rect 367336 5176 367342 5188
rect 387150 5176 387156 5188
rect 387208 5176 387214 5228
rect 412634 5176 412640 5228
rect 412692 5216 412698 5228
rect 519538 5216 519544 5228
rect 412692 5188 519544 5216
rect 412692 5176 412698 5188
rect 519538 5176 519544 5188
rect 519596 5176 519602 5228
rect 121086 5108 121092 5160
rect 121144 5148 121150 5160
rect 188338 5148 188344 5160
rect 121144 5120 188344 5148
rect 121144 5108 121150 5120
rect 188338 5108 188344 5120
rect 188396 5108 188402 5160
rect 189718 5108 189724 5160
rect 189776 5148 189782 5160
rect 299474 5148 299480 5160
rect 189776 5120 299480 5148
rect 189776 5108 189782 5120
rect 299474 5108 299480 5120
rect 299532 5108 299538 5160
rect 306742 5108 306748 5160
rect 306800 5148 306806 5160
rect 339586 5148 339592 5160
rect 306800 5120 339592 5148
rect 306800 5108 306806 5120
rect 339586 5108 339592 5120
rect 339644 5108 339650 5160
rect 371326 5108 371332 5160
rect 371384 5148 371390 5160
rect 400122 5148 400128 5160
rect 371384 5120 400128 5148
rect 371384 5108 371390 5120
rect 400122 5108 400128 5120
rect 400180 5108 400186 5160
rect 414014 5108 414020 5160
rect 414072 5148 414078 5160
rect 523034 5148 523040 5160
rect 414072 5120 523040 5148
rect 414072 5108 414078 5120
rect 523034 5108 523040 5120
rect 523092 5108 523098 5160
rect 114002 5040 114008 5092
rect 114060 5080 114066 5092
rect 181438 5080 181444 5092
rect 114060 5052 181444 5080
rect 114060 5040 114066 5052
rect 181438 5040 181444 5052
rect 181496 5040 181502 5092
rect 186130 5040 186136 5092
rect 186188 5080 186194 5092
rect 298186 5080 298192 5092
rect 186188 5052 298192 5080
rect 186188 5040 186194 5052
rect 298186 5040 298192 5052
rect 298244 5040 298250 5092
rect 303154 5040 303160 5092
rect 303212 5080 303218 5092
rect 338206 5080 338212 5092
rect 303212 5052 338212 5080
rect 303212 5040 303218 5052
rect 338206 5040 338212 5052
rect 338264 5040 338270 5092
rect 367094 5040 367100 5092
rect 367152 5080 367158 5092
rect 367278 5080 367284 5092
rect 367152 5052 367284 5080
rect 367152 5040 367158 5052
rect 367278 5040 367284 5052
rect 367336 5040 367342 5092
rect 373994 5040 374000 5092
rect 374052 5080 374058 5092
rect 407206 5080 407212 5092
rect 374052 5052 407212 5080
rect 374052 5040 374058 5052
rect 407206 5040 407212 5052
rect 407264 5040 407270 5092
rect 415394 5040 415400 5092
rect 415452 5080 415458 5092
rect 526622 5080 526628 5092
rect 415452 5052 526628 5080
rect 415452 5040 415458 5052
rect 526622 5040 526628 5052
rect 526680 5040 526686 5092
rect 103330 4972 103336 5024
rect 103388 5012 103394 5024
rect 173158 5012 173164 5024
rect 103388 4984 173164 5012
rect 103388 4972 103394 4984
rect 173158 4972 173164 4984
rect 173216 4972 173222 5024
rect 182542 4972 182548 5024
rect 182600 5012 182606 5024
rect 296806 5012 296812 5024
rect 182600 4984 296812 5012
rect 182600 4972 182606 4984
rect 296806 4972 296812 4984
rect 296864 4972 296870 5024
rect 299658 4972 299664 5024
rect 299716 5012 299722 5024
rect 336918 5012 336924 5024
rect 299716 4984 336924 5012
rect 299716 4972 299722 4984
rect 336918 4972 336924 4984
rect 336976 4972 336982 5024
rect 375374 4972 375380 5024
rect 375432 5012 375438 5024
rect 410794 5012 410800 5024
rect 375432 4984 410800 5012
rect 375432 4972 375438 4984
rect 410794 4972 410800 4984
rect 410852 4972 410858 5024
rect 416774 4972 416780 5024
rect 416832 5012 416838 5024
rect 530118 5012 530124 5024
rect 416832 4984 530124 5012
rect 416832 4972 416838 4984
rect 530118 4972 530124 4984
rect 530176 4972 530182 5024
rect 106918 4904 106924 4956
rect 106976 4944 106982 4956
rect 177298 4944 177304 4956
rect 106976 4916 177304 4944
rect 106976 4904 106982 4916
rect 177298 4904 177304 4916
rect 177356 4904 177362 4956
rect 179046 4904 179052 4956
rect 179104 4944 179110 4956
rect 295334 4944 295340 4956
rect 179104 4916 295340 4944
rect 179104 4904 179110 4916
rect 295334 4904 295340 4916
rect 295392 4904 295398 4956
rect 296070 4904 296076 4956
rect 296128 4944 296134 4956
rect 335538 4944 335544 4956
rect 296128 4916 335544 4944
rect 296128 4904 296134 4916
rect 335538 4904 335544 4916
rect 335596 4904 335602 4956
rect 376754 4904 376760 4956
rect 376812 4944 376818 4956
rect 414290 4944 414296 4956
rect 376812 4916 414296 4944
rect 376812 4904 376818 4916
rect 414290 4904 414296 4916
rect 414348 4904 414354 4956
rect 418154 4904 418160 4956
rect 418212 4944 418218 4956
rect 537202 4944 537208 4956
rect 418212 4916 537208 4944
rect 418212 4904 418218 4916
rect 537202 4904 537208 4916
rect 537260 4904 537266 4956
rect 132954 4836 132960 4888
rect 133012 4876 133018 4888
rect 280154 4876 280160 4888
rect 133012 4848 280160 4876
rect 133012 4836 133018 4848
rect 280154 4836 280160 4848
rect 280212 4836 280218 4888
rect 292574 4836 292580 4888
rect 292632 4876 292638 4888
rect 335630 4876 335636 4888
rect 292632 4848 335636 4876
rect 292632 4836 292638 4848
rect 335630 4836 335636 4848
rect 335688 4836 335694 4888
rect 378226 4836 378232 4888
rect 378284 4876 378290 4888
rect 417878 4876 417884 4888
rect 378284 4848 417884 4876
rect 378284 4836 378290 4848
rect 417878 4836 417884 4848
rect 417936 4836 417942 4888
rect 419626 4836 419632 4888
rect 419684 4876 419690 4888
rect 540790 4876 540796 4888
rect 419684 4848 540796 4876
rect 419684 4836 419690 4848
rect 540790 4836 540796 4848
rect 540848 4836 540854 4888
rect 129366 4768 129372 4820
rect 129424 4808 129430 4820
rect 278774 4808 278780 4820
rect 129424 4780 278780 4808
rect 129424 4768 129430 4780
rect 278774 4768 278780 4780
rect 278832 4768 278838 4820
rect 281902 4768 281908 4820
rect 281960 4808 281966 4820
rect 331398 4808 331404 4820
rect 281960 4780 331404 4808
rect 281960 4768 281966 4780
rect 331398 4768 331404 4780
rect 331456 4768 331462 4820
rect 378318 4768 378324 4820
rect 378376 4808 378382 4820
rect 420178 4808 420184 4820
rect 378376 4780 420184 4808
rect 378376 4768 378382 4780
rect 420178 4768 420184 4780
rect 420236 4768 420242 4820
rect 420914 4768 420920 4820
rect 420972 4808 420978 4820
rect 544378 4808 544384 4820
rect 420972 4780 544384 4808
rect 420972 4768 420978 4780
rect 544378 4768 544384 4780
rect 544436 4768 544442 4820
rect 214466 4700 214472 4752
rect 214524 4740 214530 4752
rect 307846 4740 307852 4752
rect 214524 4712 307852 4740
rect 214524 4700 214530 4712
rect 307846 4700 307852 4712
rect 307904 4700 307910 4752
rect 407114 4700 407120 4752
rect 407172 4740 407178 4752
rect 501782 4740 501788 4752
rect 407172 4712 501788 4740
rect 407172 4700 407178 4712
rect 501782 4700 501788 4712
rect 501840 4700 501846 4752
rect 218054 4632 218060 4684
rect 218112 4672 218118 4684
rect 309134 4672 309140 4684
rect 218112 4644 309140 4672
rect 218112 4632 218118 4644
rect 309134 4632 309140 4644
rect 309192 4632 309198 4684
rect 405734 4632 405740 4684
rect 405792 4672 405798 4684
rect 498194 4672 498200 4684
rect 405792 4644 498200 4672
rect 405792 4632 405798 4644
rect 498194 4632 498200 4644
rect 498252 4632 498258 4684
rect 175458 4564 175464 4616
rect 175516 4604 175522 4616
rect 260098 4604 260104 4616
rect 175516 4576 260104 4604
rect 175516 4564 175522 4576
rect 260098 4564 260104 4576
rect 260156 4564 260162 4616
rect 299290 4564 299296 4616
rect 299348 4604 299354 4616
rect 329834 4604 329840 4616
rect 299348 4576 329840 4604
rect 299348 4564 299354 4576
rect 329834 4564 329840 4576
rect 329892 4564 329898 4616
rect 379606 4564 379612 4616
rect 379664 4604 379670 4616
rect 423766 4604 423772 4616
rect 379664 4576 423772 4604
rect 379664 4564 379670 4576
rect 423766 4564 423772 4576
rect 423824 4564 423830 4616
rect 298002 4496 298008 4548
rect 298060 4536 298066 4548
rect 324314 4536 324320 4548
rect 298060 4508 324320 4536
rect 298060 4496 298066 4508
rect 324314 4496 324320 4508
rect 324372 4496 324378 4548
rect 379514 4496 379520 4548
rect 379572 4536 379578 4548
rect 421374 4536 421380 4548
rect 379572 4508 421380 4536
rect 379572 4496 379578 4508
rect 421374 4496 421380 4508
rect 421432 4496 421438 4548
rect 299382 4428 299388 4480
rect 299440 4468 299446 4480
rect 324222 4468 324228 4480
rect 299440 4440 324228 4468
rect 299440 4428 299446 4440
rect 324222 4428 324228 4440
rect 324280 4428 324286 4480
rect 378134 4428 378140 4480
rect 378192 4468 378198 4480
rect 418982 4468 418988 4480
rect 378192 4440 418988 4468
rect 378192 4428 378198 4440
rect 418982 4428 418988 4440
rect 419040 4428 419046 4480
rect 301498 4360 301504 4412
rect 301556 4400 301562 4412
rect 325786 4400 325792 4412
rect 301556 4372 325792 4400
rect 301556 4360 301562 4372
rect 325786 4360 325792 4372
rect 325844 4360 325850 4412
rect 328730 4332 328736 4344
rect 306346 4304 328736 4332
rect 306346 4264 306374 4304
rect 328730 4292 328736 4304
rect 328788 4292 328794 4344
rect 303632 4236 306374 4264
rect 176654 4156 176660 4208
rect 176712 4196 176718 4208
rect 177850 4196 177856 4208
rect 176712 4168 177856 4196
rect 176712 4156 176718 4168
rect 177850 4156 177856 4168
rect 177908 4156 177914 4208
rect 226334 4156 226340 4208
rect 226392 4196 226398 4208
rect 227530 4196 227536 4208
rect 226392 4168 227536 4196
rect 226392 4156 226398 4168
rect 227530 4156 227536 4168
rect 227588 4156 227594 4208
rect 99834 4088 99840 4140
rect 99892 4128 99898 4140
rect 269206 4128 269212 4140
rect 99892 4100 269212 4128
rect 99892 4088 99898 4100
rect 269206 4088 269212 4100
rect 269264 4088 269270 4140
rect 274818 4088 274824 4140
rect 274876 4128 274882 4140
rect 303632 4128 303660 4236
rect 378888 4168 379100 4196
rect 274876 4100 303660 4128
rect 274876 4088 274882 4100
rect 311434 4088 311440 4140
rect 311492 4128 311498 4140
rect 340874 4128 340880 4140
rect 311492 4100 340880 4128
rect 311492 4088 311498 4100
rect 340874 4088 340880 4100
rect 340932 4088 340938 4140
rect 342162 4088 342168 4140
rect 342220 4128 342226 4140
rect 352098 4128 352104 4140
rect 342220 4100 352104 4128
rect 342220 4088 342226 4100
rect 352098 4088 352104 4100
rect 352156 4088 352162 4140
rect 363230 4088 363236 4140
rect 363288 4128 363294 4140
rect 367094 4128 367100 4140
rect 363288 4100 367100 4128
rect 363288 4088 363294 4100
rect 367094 4088 367100 4100
rect 367152 4088 367158 4140
rect 367186 4088 367192 4140
rect 367244 4128 367250 4140
rect 378778 4128 378784 4140
rect 367244 4100 378784 4128
rect 367244 4088 367250 4100
rect 378778 4088 378784 4100
rect 378836 4088 378842 4140
rect 92750 4020 92756 4072
rect 92808 4060 92814 4072
rect 266446 4060 266452 4072
rect 92808 4032 266452 4060
rect 92808 4020 92814 4032
rect 266446 4020 266452 4032
rect 266504 4020 266510 4072
rect 267734 4020 267740 4072
rect 267792 4060 267798 4072
rect 301498 4060 301504 4072
rect 267792 4032 301504 4060
rect 267792 4020 267798 4032
rect 301498 4020 301504 4032
rect 301556 4020 301562 4072
rect 309042 4020 309048 4072
rect 309100 4060 309106 4072
rect 340782 4060 340788 4072
rect 309100 4032 340788 4060
rect 309100 4020 309106 4032
rect 340782 4020 340788 4032
rect 340840 4020 340846 4072
rect 340966 4020 340972 4072
rect 341024 4060 341030 4072
rect 341024 4032 350856 4060
rect 341024 4020 341030 4032
rect 82078 3952 82084 4004
rect 82136 3992 82142 4004
rect 262214 3992 262220 4004
rect 82136 3964 262220 3992
rect 82136 3952 82142 3964
rect 262214 3952 262220 3964
rect 262272 3952 262278 4004
rect 264146 3952 264152 4004
rect 264204 3992 264210 4004
rect 299382 3992 299388 4004
rect 264204 3964 299388 3992
rect 264204 3952 264210 3964
rect 299382 3952 299388 3964
rect 299440 3952 299446 4004
rect 317874 3952 317880 4004
rect 317932 3992 317938 4004
rect 322934 3992 322940 4004
rect 317932 3964 322940 3992
rect 317932 3952 317938 3964
rect 322934 3952 322940 3964
rect 322992 3952 322998 4004
rect 338666 3952 338672 4004
rect 338724 3992 338730 4004
rect 350718 3992 350724 4004
rect 338724 3964 350724 3992
rect 338724 3952 338730 3964
rect 350718 3952 350724 3964
rect 350776 3952 350782 4004
rect 350828 3992 350856 4032
rect 351638 4020 351644 4072
rect 351696 4060 351702 4072
rect 354766 4060 354772 4072
rect 351696 4032 354772 4060
rect 351696 4020 351702 4032
rect 354766 4020 354772 4032
rect 354824 4020 354830 4072
rect 360838 4020 360844 4072
rect 360896 4060 360902 4072
rect 364610 4060 364616 4072
rect 360896 4032 364616 4060
rect 360896 4020 360902 4032
rect 364610 4020 364616 4032
rect 364668 4020 364674 4072
rect 365714 4020 365720 4072
rect 365772 4060 365778 4072
rect 378888 4060 378916 4168
rect 379072 4128 379100 4168
rect 400858 4156 400864 4208
rect 400916 4196 400922 4208
rect 400916 4168 402652 4196
rect 400916 4156 400922 4168
rect 379072 4100 379514 4128
rect 365772 4032 378916 4060
rect 379486 4060 379514 4100
rect 383654 4088 383660 4140
rect 383712 4128 383718 4140
rect 383712 4100 384896 4128
rect 383712 4088 383718 4100
rect 384758 4060 384764 4072
rect 379486 4032 384764 4060
rect 365772 4020 365778 4032
rect 384758 4020 384764 4032
rect 384816 4020 384822 4072
rect 384868 4060 384896 4100
rect 388346 4088 388352 4140
rect 388404 4128 388410 4140
rect 402514 4128 402520 4140
rect 388404 4100 402520 4128
rect 388404 4088 388410 4100
rect 402514 4088 402520 4100
rect 402572 4088 402578 4140
rect 402624 4128 402652 4168
rect 403618 4128 403624 4140
rect 402624 4100 403624 4128
rect 403618 4088 403624 4100
rect 403676 4088 403682 4140
rect 404998 4088 405004 4140
rect 405056 4128 405062 4140
rect 411898 4128 411904 4140
rect 405056 4100 411904 4128
rect 405056 4088 405062 4100
rect 411898 4088 411904 4100
rect 411956 4088 411962 4140
rect 411990 4088 411996 4140
rect 412048 4128 412054 4140
rect 440326 4128 440332 4140
rect 412048 4100 440332 4128
rect 412048 4088 412054 4100
rect 440326 4088 440332 4100
rect 440384 4088 440390 4140
rect 440970 4088 440976 4140
rect 441028 4128 441034 4140
rect 550266 4128 550272 4140
rect 441028 4100 550272 4128
rect 441028 4088 441034 4100
rect 550266 4088 550272 4100
rect 550324 4088 550330 4140
rect 384868 4032 388392 4060
rect 352190 3992 352196 4004
rect 350828 3964 352196 3992
rect 352190 3952 352196 3964
rect 352248 3952 352254 4004
rect 360286 3952 360292 4004
rect 360344 3992 360350 4004
rect 367002 3992 367008 4004
rect 360344 3964 367008 3992
rect 360344 3952 360350 3964
rect 367002 3952 367008 3964
rect 367060 3952 367066 4004
rect 368474 3952 368480 4004
rect 368532 3992 368538 4004
rect 368532 3964 372844 3992
rect 368532 3952 368538 3964
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 248690 3924 248696 3936
rect 43128 3896 248696 3924
rect 43128 3884 43134 3896
rect 248690 3884 248696 3896
rect 248748 3884 248754 3936
rect 276014 3884 276020 3936
rect 276072 3924 276078 3936
rect 288526 3924 288532 3936
rect 276072 3896 288532 3924
rect 276072 3884 276078 3896
rect 288526 3884 288532 3896
rect 288584 3884 288590 3936
rect 294874 3884 294880 3936
rect 294932 3924 294938 3936
rect 335354 3924 335360 3936
rect 294932 3896 335360 3924
rect 294932 3884 294938 3896
rect 335354 3884 335360 3896
rect 335412 3884 335418 3936
rect 336274 3884 336280 3936
rect 336332 3924 336338 3936
rect 349246 3924 349252 3936
rect 336332 3896 349252 3924
rect 336332 3884 336338 3896
rect 349246 3884 349252 3896
rect 349304 3884 349310 3936
rect 363138 3884 363144 3936
rect 363196 3924 363202 3936
rect 372816 3924 372844 3964
rect 377398 3952 377404 4004
rect 377456 3992 377462 4004
rect 378870 3992 378876 4004
rect 377456 3964 378876 3992
rect 377456 3952 377462 3964
rect 378870 3952 378876 3964
rect 378928 3952 378934 4004
rect 378962 3952 378968 4004
rect 379020 3992 379026 4004
rect 388254 3992 388260 4004
rect 379020 3964 388260 3992
rect 379020 3952 379026 3964
rect 388254 3952 388260 3964
rect 388312 3952 388318 4004
rect 388364 3992 388392 4032
rect 391198 4020 391204 4072
rect 391256 4060 391262 4072
rect 413094 4060 413100 4072
rect 391256 4032 413100 4060
rect 391256 4020 391262 4032
rect 413094 4020 413100 4032
rect 413152 4020 413158 4072
rect 416038 4020 416044 4072
rect 416096 4060 416102 4072
rect 447410 4060 447416 4072
rect 416096 4032 447416 4060
rect 416096 4020 416102 4032
rect 447410 4020 447416 4032
rect 447468 4020 447474 4072
rect 447778 4020 447784 4072
rect 447836 4060 447842 4072
rect 557350 4060 557356 4072
rect 447836 4032 557356 4060
rect 447836 4020 447842 4032
rect 557350 4020 557356 4032
rect 557408 4020 557414 4072
rect 393130 3992 393136 4004
rect 388364 3964 393136 3992
rect 393130 3952 393136 3964
rect 393188 3952 393194 4004
rect 402698 3952 402704 4004
rect 402756 3992 402762 4004
rect 404814 3992 404820 4004
rect 402756 3964 404820 3992
rect 402756 3952 402762 3964
rect 404814 3952 404820 3964
rect 404872 3952 404878 4004
rect 405734 3952 405740 4004
rect 405792 3992 405798 4004
rect 472250 3992 472256 4004
rect 405792 3964 472256 3992
rect 405792 3952 405798 3964
rect 472250 3952 472256 3964
rect 472308 3952 472314 4004
rect 472618 3952 472624 4004
rect 472676 3992 472682 4004
rect 582190 3992 582196 4004
rect 472676 3964 582196 3992
rect 472676 3952 472682 3964
rect 582190 3952 582196 3964
rect 582248 3952 582254 4004
rect 363196 3896 371004 3924
rect 372816 3896 379514 3924
rect 363196 3884 363202 3896
rect 35986 3816 35992 3868
rect 36044 3856 36050 3868
rect 247034 3856 247040 3868
rect 36044 3828 247040 3856
rect 36044 3816 36050 3828
rect 247034 3816 247040 3828
rect 247092 3816 247098 3868
rect 248782 3816 248788 3868
rect 248840 3856 248846 3868
rect 290734 3856 290740 3868
rect 248840 3828 290740 3856
rect 248840 3816 248846 3828
rect 290734 3816 290740 3828
rect 290792 3816 290798 3868
rect 293678 3816 293684 3868
rect 293736 3856 293742 3868
rect 335446 3856 335452 3868
rect 293736 3828 335452 3856
rect 293736 3816 293742 3828
rect 335446 3816 335452 3828
rect 335504 3816 335510 3868
rect 337470 3816 337476 3868
rect 337528 3856 337534 3868
rect 350626 3856 350632 3868
rect 337528 3828 350632 3856
rect 337528 3816 337534 3828
rect 350626 3816 350632 3828
rect 350684 3816 350690 3868
rect 363046 3816 363052 3868
rect 363104 3856 363110 3868
rect 370866 3856 370872 3868
rect 363104 3828 370872 3856
rect 363104 3816 363110 3828
rect 370866 3816 370872 3828
rect 370924 3816 370930 3868
rect 370976 3856 371004 3896
rect 374086 3856 374092 3868
rect 370976 3828 374092 3856
rect 374086 3816 374092 3828
rect 374144 3816 374150 3868
rect 379486 3856 379514 3896
rect 382274 3884 382280 3936
rect 382332 3924 382338 3936
rect 433242 3924 433248 3936
rect 382332 3896 433248 3924
rect 382332 3884 382338 3896
rect 433242 3884 433248 3896
rect 433300 3884 433306 3936
rect 433886 3884 433892 3936
rect 433944 3924 433950 3936
rect 450906 3924 450912 3936
rect 433944 3896 450912 3924
rect 433944 3884 433950 3896
rect 450906 3884 450912 3896
rect 450964 3884 450970 3936
rect 451918 3884 451924 3936
rect 451976 3924 451982 3936
rect 564434 3924 564440 3936
rect 451976 3896 564440 3924
rect 451976 3884 451982 3896
rect 564434 3884 564440 3896
rect 564492 3884 564498 3936
rect 390646 3856 390652 3868
rect 379486 3828 390652 3856
rect 390646 3816 390652 3828
rect 390704 3816 390710 3868
rect 391934 3816 391940 3868
rect 391992 3856 391998 3868
rect 458082 3856 458088 3868
rect 391992 3828 458088 3856
rect 391992 3816 391998 3828
rect 458082 3816 458088 3828
rect 458140 3816 458146 3868
rect 458818 3816 458824 3868
rect 458876 3856 458882 3868
rect 578602 3856 578608 3868
rect 458876 3828 578608 3856
rect 458876 3816 458882 3828
rect 578602 3816 578608 3828
rect 578660 3816 578666 3868
rect 28902 3748 28908 3800
rect 28960 3788 28966 3800
rect 244274 3788 244280 3800
rect 28960 3760 244280 3788
rect 28960 3748 28966 3760
rect 244274 3748 244280 3760
rect 244332 3748 244338 3800
rect 245194 3748 245200 3800
rect 245252 3788 245258 3800
rect 264238 3788 264244 3800
rect 245252 3760 264244 3788
rect 245252 3748 245258 3760
rect 264238 3748 264244 3760
rect 264296 3748 264302 3800
rect 280706 3748 280712 3800
rect 280764 3788 280770 3800
rect 331306 3788 331312 3800
rect 280764 3760 331312 3788
rect 280764 3748 280770 3760
rect 331306 3748 331312 3760
rect 331364 3748 331370 3800
rect 332686 3748 332692 3800
rect 332744 3788 332750 3800
rect 349522 3788 349528 3800
rect 332744 3760 349528 3788
rect 332744 3748 332750 3760
rect 349522 3748 349528 3760
rect 349580 3748 349586 3800
rect 363322 3748 363328 3800
rect 363380 3788 363386 3800
rect 363690 3788 363696 3800
rect 363380 3760 363696 3788
rect 363380 3748 363386 3760
rect 363690 3748 363696 3760
rect 363748 3748 363754 3800
rect 367094 3748 367100 3800
rect 367152 3788 367158 3800
rect 375282 3788 375288 3800
rect 367152 3760 375288 3788
rect 367152 3748 367158 3760
rect 375282 3748 375288 3760
rect 375340 3748 375346 3800
rect 376018 3748 376024 3800
rect 376076 3788 376082 3800
rect 398926 3788 398932 3800
rect 376076 3760 398932 3788
rect 376076 3748 376082 3760
rect 398926 3748 398932 3760
rect 398984 3748 398990 3800
rect 402606 3748 402612 3800
rect 402664 3788 402670 3800
rect 408402 3788 408408 3800
rect 402664 3760 408408 3788
rect 402664 3748 402670 3760
rect 408402 3748 408408 3760
rect 408460 3748 408466 3800
rect 409138 3748 409144 3800
rect 409196 3788 409202 3800
rect 415486 3788 415492 3800
rect 409196 3760 415492 3788
rect 409196 3748 409202 3760
rect 415486 3748 415492 3760
rect 415544 3748 415550 3800
rect 419534 3748 419540 3800
rect 419592 3788 419598 3800
rect 539594 3788 539600 3800
rect 419592 3760 539600 3788
rect 419592 3748 419598 3760
rect 539594 3748 539600 3760
rect 539652 3748 539658 3800
rect 24210 3680 24216 3732
rect 24268 3720 24274 3732
rect 243078 3720 243084 3732
rect 24268 3692 243084 3720
rect 24268 3680 24274 3692
rect 243078 3680 243084 3692
rect 243136 3680 243142 3732
rect 257062 3680 257068 3732
rect 257120 3720 257126 3732
rect 317874 3720 317880 3732
rect 257120 3692 317880 3720
rect 257120 3680 257126 3692
rect 317874 3680 317880 3692
rect 317932 3680 317938 3732
rect 321554 3720 321560 3732
rect 317984 3692 321560 3720
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 241606 3652 241612 3664
rect 20680 3624 241612 3652
rect 20680 3612 20686 3624
rect 241606 3612 241612 3624
rect 241664 3612 241670 3664
rect 253474 3612 253480 3664
rect 253532 3652 253538 3664
rect 317984 3652 318012 3692
rect 321554 3680 321560 3692
rect 321612 3680 321618 3732
rect 330386 3680 330392 3732
rect 330444 3720 330450 3732
rect 347866 3720 347872 3732
rect 330444 3692 347872 3720
rect 330444 3680 330450 3692
rect 347866 3680 347872 3692
rect 347924 3680 347930 3732
rect 360194 3680 360200 3732
rect 360252 3720 360258 3732
rect 360252 3692 364334 3720
rect 360252 3680 360258 3692
rect 320174 3652 320180 3664
rect 253532 3624 318012 3652
rect 318076 3624 320180 3652
rect 253532 3612 253538 3624
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 241514 3584 241520 3596
rect 19484 3556 241520 3584
rect 19484 3544 19490 3556
rect 241514 3544 241520 3556
rect 241572 3544 241578 3596
rect 249978 3544 249984 3596
rect 250036 3584 250042 3596
rect 318076 3584 318104 3624
rect 320174 3612 320180 3624
rect 320232 3612 320238 3664
rect 325602 3612 325608 3664
rect 325660 3652 325666 3664
rect 346486 3652 346492 3664
rect 325660 3624 346492 3652
rect 325660 3612 325666 3624
rect 346486 3612 346492 3624
rect 346544 3612 346550 3664
rect 349246 3612 349252 3664
rect 349304 3652 349310 3664
rect 354858 3652 354864 3664
rect 349304 3624 354864 3652
rect 349304 3612 349310 3624
rect 354858 3612 354864 3624
rect 354916 3612 354922 3664
rect 361574 3612 361580 3664
rect 361632 3652 361638 3664
rect 364306 3652 364334 3692
rect 365806 3680 365812 3732
rect 365864 3720 365870 3732
rect 381170 3720 381176 3732
rect 365864 3692 381176 3720
rect 365864 3680 365870 3692
rect 381170 3680 381176 3692
rect 381228 3680 381234 3732
rect 388438 3680 388444 3732
rect 388496 3720 388502 3732
rect 393038 3720 393044 3732
rect 388496 3692 393044 3720
rect 388496 3680 388502 3692
rect 393038 3680 393044 3692
rect 393096 3680 393102 3732
rect 393130 3680 393136 3732
rect 393188 3720 393194 3732
rect 436738 3720 436744 3732
rect 393188 3692 436744 3720
rect 393188 3680 393194 3692
rect 436738 3680 436744 3692
rect 436796 3680 436802 3732
rect 450538 3680 450544 3732
rect 450596 3720 450602 3732
rect 571518 3720 571524 3732
rect 450596 3692 571524 3720
rect 450596 3680 450602 3692
rect 571518 3680 571524 3692
rect 571576 3680 571582 3732
rect 368198 3652 368204 3664
rect 361632 3624 363460 3652
rect 364306 3624 368204 3652
rect 361632 3612 361638 3624
rect 250036 3556 318104 3584
rect 250036 3544 250042 3556
rect 318886 3544 318892 3596
rect 318944 3544 318950 3596
rect 323302 3544 323308 3596
rect 323360 3584 323366 3596
rect 345198 3584 345204 3596
rect 323360 3556 345204 3584
rect 323360 3544 323366 3556
rect 345198 3544 345204 3556
rect 345256 3544 345262 3596
rect 363432 3584 363460 3624
rect 368198 3612 368204 3624
rect 368256 3612 368262 3664
rect 370866 3612 370872 3664
rect 370924 3652 370930 3664
rect 376478 3652 376484 3664
rect 370924 3624 376484 3652
rect 370924 3612 370930 3624
rect 376478 3612 376484 3624
rect 376536 3612 376542 3664
rect 376570 3612 376576 3664
rect 376628 3652 376634 3664
rect 394234 3652 394240 3664
rect 376628 3624 394240 3652
rect 376628 3612 376634 3624
rect 394234 3612 394240 3624
rect 394292 3612 394298 3664
rect 394326 3612 394332 3664
rect 394384 3652 394390 3664
rect 401318 3652 401324 3664
rect 394384 3624 401324 3652
rect 394384 3612 394390 3624
rect 401318 3612 401324 3624
rect 401376 3612 401382 3664
rect 406378 3612 406384 3664
rect 406436 3652 406442 3664
rect 406436 3624 412036 3652
rect 406436 3612 406442 3624
rect 369394 3584 369400 3596
rect 363432 3556 369400 3584
rect 369394 3544 369400 3556
rect 369452 3544 369458 3596
rect 371234 3544 371240 3596
rect 371292 3584 371298 3596
rect 397730 3584 397736 3596
rect 371292 3556 397736 3584
rect 371292 3544 371298 3556
rect 397730 3544 397736 3556
rect 397788 3544 397794 3596
rect 398098 3544 398104 3596
rect 398156 3584 398162 3596
rect 402698 3584 402704 3596
rect 398156 3556 402704 3584
rect 398156 3544 398162 3556
rect 402698 3544 402704 3556
rect 402756 3544 402762 3596
rect 406470 3544 406476 3596
rect 406528 3584 406534 3596
rect 411898 3584 411904 3596
rect 406528 3556 411904 3584
rect 406528 3544 406534 3556
rect 411898 3544 411904 3556
rect 411956 3544 411962 3596
rect 412008 3584 412036 3624
rect 412082 3612 412088 3664
rect 412140 3652 412146 3664
rect 416682 3652 416688 3664
rect 412140 3624 416688 3652
rect 412140 3612 412146 3624
rect 416682 3612 416688 3624
rect 416740 3612 416746 3664
rect 423674 3612 423680 3664
rect 423732 3652 423738 3664
rect 553762 3652 553768 3664
rect 423732 3624 553768 3652
rect 423732 3612 423738 3624
rect 553762 3612 553768 3624
rect 553820 3612 553826 3664
rect 422570 3584 422576 3596
rect 412008 3556 422576 3584
rect 422570 3544 422576 3556
rect 422628 3544 422634 3596
rect 426434 3544 426440 3596
rect 426492 3584 426498 3596
rect 560846 3584 560852 3596
rect 426492 3556 560852 3584
rect 426492 3544 426498 3556
rect 560846 3544 560852 3556
rect 560904 3544 560910 3596
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 238754 3516 238760 3528
rect 14792 3488 238760 3516
rect 14792 3476 14798 3488
rect 238754 3476 238760 3488
rect 238812 3476 238818 3528
rect 246390 3476 246396 3528
rect 246448 3516 246454 3528
rect 318904 3516 318932 3544
rect 246448 3488 318932 3516
rect 246448 3476 246454 3488
rect 322106 3476 322112 3528
rect 322164 3516 322170 3528
rect 345106 3516 345112 3528
rect 322164 3488 345112 3516
rect 322164 3476 322170 3488
rect 345106 3476 345112 3488
rect 345164 3476 345170 3528
rect 352006 3516 352012 3528
rect 345492 3488 352012 3516
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 238846 3448 238852 3460
rect 11204 3420 238852 3448
rect 11204 3408 11210 3420
rect 238846 3408 238852 3420
rect 238904 3408 238910 3460
rect 242894 3408 242900 3460
rect 242952 3448 242958 3460
rect 317414 3448 317420 3460
rect 242952 3420 317420 3448
rect 242952 3408 242958 3420
rect 317414 3408 317420 3420
rect 317472 3408 317478 3460
rect 329190 3408 329196 3460
rect 329248 3448 329254 3460
rect 333238 3448 333244 3460
rect 329248 3420 333244 3448
rect 329248 3408 329254 3420
rect 333238 3408 333244 3420
rect 333296 3408 333302 3460
rect 333882 3408 333888 3460
rect 333940 3448 333946 3460
rect 334618 3448 334624 3460
rect 333940 3420 334624 3448
rect 333940 3408 333946 3420
rect 334618 3408 334624 3420
rect 334676 3408 334682 3460
rect 344554 3408 344560 3460
rect 344612 3448 344618 3460
rect 345492 3448 345520 3488
rect 352006 3476 352012 3488
rect 352064 3476 352070 3528
rect 352834 3476 352840 3528
rect 352892 3516 352898 3528
rect 353938 3516 353944 3528
rect 352892 3488 353944 3516
rect 352892 3476 352898 3488
rect 353938 3476 353944 3488
rect 353996 3476 354002 3528
rect 355226 3476 355232 3528
rect 355284 3516 355290 3528
rect 356238 3516 356244 3528
rect 355284 3488 356244 3516
rect 355284 3476 355290 3488
rect 356238 3476 356244 3488
rect 356296 3476 356302 3528
rect 357526 3476 357532 3528
rect 357584 3516 357590 3528
rect 358722 3516 358728 3528
rect 357584 3488 358728 3516
rect 357584 3476 357590 3488
rect 358722 3476 358728 3488
rect 358780 3476 358786 3528
rect 358906 3476 358912 3528
rect 358964 3516 358970 3528
rect 361114 3516 361120 3528
rect 358964 3488 361120 3516
rect 358964 3476 358970 3488
rect 361114 3476 361120 3488
rect 361172 3476 361178 3528
rect 364334 3476 364340 3528
rect 364392 3516 364398 3528
rect 377674 3516 377680 3528
rect 364392 3488 377680 3516
rect 364392 3476 364398 3488
rect 377674 3476 377680 3488
rect 377732 3476 377738 3528
rect 380250 3476 380256 3528
rect 380308 3516 380314 3528
rect 388346 3516 388352 3528
rect 380308 3488 388352 3516
rect 380308 3476 380314 3488
rect 388346 3476 388352 3488
rect 388404 3476 388410 3528
rect 388438 3476 388444 3528
rect 388496 3516 388502 3528
rect 426158 3516 426164 3528
rect 388496 3488 426164 3516
rect 388496 3476 388502 3488
rect 426158 3476 426164 3488
rect 426216 3476 426222 3528
rect 431954 3476 431960 3528
rect 432012 3516 432018 3528
rect 575106 3516 575112 3528
rect 432012 3488 575112 3516
rect 432012 3476 432018 3488
rect 575106 3476 575112 3488
rect 575164 3476 575170 3528
rect 349338 3448 349344 3460
rect 344612 3420 345520 3448
rect 345584 3420 349344 3448
rect 344612 3408 344618 3420
rect 44174 3340 44180 3392
rect 44232 3380 44238 3392
rect 45094 3380 45100 3392
rect 44232 3352 45100 3380
rect 44232 3340 44238 3352
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 52454 3340 52460 3392
rect 52512 3380 52518 3392
rect 53374 3380 53380 3392
rect 52512 3352 53380 3380
rect 52512 3340 52518 3352
rect 53374 3340 53380 3352
rect 53432 3340 53438 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 271874 3380 271880 3392
rect 113146 3352 271880 3380
rect 110506 3272 110512 3324
rect 110564 3312 110570 3324
rect 113146 3312 113174 3352
rect 271874 3340 271880 3352
rect 271932 3340 271938 3392
rect 278314 3340 278320 3392
rect 278372 3380 278378 3392
rect 299290 3380 299296 3392
rect 278372 3352 299296 3380
rect 278372 3340 278378 3352
rect 299290 3340 299296 3352
rect 299348 3340 299354 3392
rect 315022 3340 315028 3392
rect 315080 3380 315086 3392
rect 342438 3380 342444 3392
rect 315080 3352 342444 3380
rect 315080 3340 315086 3352
rect 342438 3340 342444 3352
rect 342496 3340 342502 3392
rect 110564 3284 113174 3312
rect 110564 3272 110570 3284
rect 117590 3272 117596 3324
rect 117648 3312 117654 3324
rect 274634 3312 274640 3324
rect 117648 3284 274640 3312
rect 117648 3272 117654 3284
rect 274634 3272 274640 3284
rect 274692 3272 274698 3324
rect 300762 3272 300768 3324
rect 300820 3312 300826 3324
rect 326430 3312 326436 3324
rect 300820 3284 326436 3312
rect 300820 3272 300826 3284
rect 326430 3272 326436 3284
rect 326488 3272 326494 3324
rect 335078 3272 335084 3324
rect 335136 3312 335142 3324
rect 345584 3312 345612 3420
rect 349338 3408 349344 3420
rect 349396 3408 349402 3460
rect 364426 3408 364432 3460
rect 364484 3448 364490 3460
rect 364484 3420 379514 3448
rect 364484 3408 364490 3420
rect 348050 3340 348056 3392
rect 348108 3380 348114 3392
rect 353478 3380 353484 3392
rect 348108 3352 353484 3380
rect 348108 3340 348114 3352
rect 353478 3340 353484 3352
rect 353536 3340 353542 3392
rect 361666 3340 361672 3392
rect 361724 3380 361730 3392
rect 371694 3380 371700 3392
rect 361724 3352 371700 3380
rect 361724 3340 361730 3352
rect 371694 3340 371700 3352
rect 371752 3340 371758 3392
rect 379486 3380 379514 3420
rect 382366 3408 382372 3460
rect 382424 3448 382430 3460
rect 429654 3448 429660 3460
rect 382424 3420 429660 3448
rect 382424 3408 382430 3420
rect 429654 3408 429660 3420
rect 429712 3408 429718 3460
rect 433334 3408 433340 3460
rect 433392 3448 433398 3460
rect 580994 3448 581000 3460
rect 433392 3420 581000 3448
rect 433392 3408 433398 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 379974 3380 379980 3392
rect 379486 3352 379980 3380
rect 379974 3340 379980 3352
rect 380032 3340 380038 3392
rect 380066 3340 380072 3392
rect 380124 3380 380130 3392
rect 395338 3380 395344 3392
rect 380124 3352 395344 3380
rect 380124 3340 380130 3352
rect 395338 3340 395344 3352
rect 395396 3340 395402 3392
rect 396166 3340 396172 3392
rect 396224 3380 396230 3392
rect 405734 3380 405740 3392
rect 396224 3352 405740 3380
rect 396224 3340 396230 3352
rect 405734 3340 405740 3352
rect 405792 3340 405798 3392
rect 440878 3340 440884 3392
rect 440936 3380 440942 3392
rect 543182 3380 543188 3392
rect 440936 3352 543188 3380
rect 440936 3340 440942 3352
rect 543182 3340 543188 3352
rect 543240 3340 543246 3392
rect 335136 3284 345612 3312
rect 335136 3272 335142 3284
rect 346946 3272 346952 3324
rect 347004 3312 347010 3324
rect 353386 3312 353392 3324
rect 347004 3284 353392 3312
rect 347004 3272 347010 3284
rect 353386 3272 353392 3284
rect 353444 3272 353450 3324
rect 354030 3272 354036 3324
rect 354088 3312 354094 3324
rect 356146 3312 356152 3324
rect 354088 3284 356152 3312
rect 354088 3272 354094 3284
rect 356146 3272 356152 3284
rect 356204 3272 356210 3324
rect 367278 3272 367284 3324
rect 367336 3312 367342 3324
rect 385954 3312 385960 3324
rect 367336 3284 385960 3312
rect 367336 3272 367342 3284
rect 385954 3272 385960 3284
rect 386012 3272 386018 3324
rect 387058 3272 387064 3324
rect 387116 3312 387122 3324
rect 387116 3284 393314 3312
rect 387116 3272 387122 3284
rect 124674 3204 124680 3256
rect 124732 3244 124738 3256
rect 236638 3244 236644 3256
rect 124732 3216 236644 3244
rect 124732 3204 124738 3216
rect 236638 3204 236644 3216
rect 236696 3204 236702 3256
rect 260650 3204 260656 3256
rect 260708 3244 260714 3256
rect 298002 3244 298008 3256
rect 260708 3216 298008 3244
rect 260708 3204 260714 3216
rect 298002 3204 298008 3216
rect 298060 3204 298066 3256
rect 304350 3204 304356 3256
rect 304408 3244 304414 3256
rect 329098 3244 329104 3256
rect 304408 3216 329104 3244
rect 304408 3204 304414 3216
rect 329098 3204 329104 3216
rect 329156 3204 329162 3256
rect 339862 3204 339868 3256
rect 339920 3244 339926 3256
rect 350534 3244 350540 3256
rect 339920 3216 350540 3244
rect 339920 3204 339926 3216
rect 350534 3204 350540 3216
rect 350592 3204 350598 3256
rect 363690 3204 363696 3256
rect 363748 3244 363754 3256
rect 372890 3244 372896 3256
rect 363748 3216 372896 3244
rect 363748 3204 363754 3216
rect 372890 3204 372896 3216
rect 372948 3204 372954 3256
rect 374730 3204 374736 3256
rect 374788 3244 374794 3256
rect 383562 3244 383568 3256
rect 374788 3216 383568 3244
rect 374788 3204 374794 3216
rect 383562 3204 383568 3216
rect 383620 3204 383626 3256
rect 384298 3204 384304 3256
rect 384356 3244 384362 3256
rect 389450 3244 389456 3256
rect 384356 3216 389456 3244
rect 384356 3204 384362 3216
rect 389450 3204 389456 3216
rect 389508 3204 389514 3256
rect 393286 3244 393314 3284
rect 397454 3272 397460 3324
rect 397512 3312 397518 3324
rect 475746 3312 475752 3324
rect 397512 3284 475752 3312
rect 397512 3272 397518 3284
rect 475746 3272 475752 3284
rect 475804 3272 475810 3324
rect 558546 3312 558552 3324
rect 480226 3284 558552 3312
rect 406010 3244 406016 3256
rect 393286 3216 406016 3244
rect 406010 3204 406016 3216
rect 406068 3204 406074 3256
rect 460198 3204 460204 3256
rect 460256 3244 460262 3256
rect 465166 3244 465172 3256
rect 460256 3216 465172 3244
rect 460256 3204 460262 3216
rect 465166 3204 465172 3216
rect 465224 3204 465230 3256
rect 475378 3204 475384 3256
rect 475436 3244 475442 3256
rect 480226 3244 480254 3284
rect 558546 3272 558552 3284
rect 558604 3272 558610 3324
rect 475436 3216 480254 3244
rect 475436 3204 475442 3216
rect 247586 3136 247592 3188
rect 247644 3176 247650 3188
rect 261478 3176 261484 3188
rect 247644 3148 261484 3176
rect 247644 3136 247650 3148
rect 261478 3136 261484 3148
rect 261536 3136 261542 3188
rect 290182 3136 290188 3188
rect 290240 3176 290246 3188
rect 309870 3176 309876 3188
rect 290240 3148 309876 3176
rect 290240 3136 290246 3148
rect 309870 3136 309876 3148
rect 309928 3136 309934 3188
rect 320910 3136 320916 3188
rect 320968 3176 320974 3188
rect 331858 3176 331864 3188
rect 320968 3148 331864 3176
rect 320968 3136 320974 3148
rect 331858 3136 331864 3148
rect 331916 3136 331922 3188
rect 343358 3136 343364 3188
rect 343416 3176 343422 3188
rect 351914 3176 351920 3188
rect 343416 3148 351920 3176
rect 343416 3136 343422 3148
rect 351914 3136 351920 3148
rect 351972 3136 351978 3188
rect 358998 3136 359004 3188
rect 359056 3176 359062 3188
rect 362310 3176 362316 3188
rect 359056 3148 362316 3176
rect 359056 3136 359062 3148
rect 362310 3136 362316 3148
rect 362368 3136 362374 3188
rect 363598 3136 363604 3188
rect 363656 3176 363662 3188
rect 370590 3176 370596 3188
rect 363656 3148 370596 3176
rect 363656 3136 363662 3148
rect 370590 3136 370596 3148
rect 370648 3136 370654 3188
rect 374638 3136 374644 3188
rect 374696 3176 374702 3188
rect 380066 3176 380072 3188
rect 374696 3148 380072 3176
rect 374696 3136 374702 3148
rect 380066 3136 380072 3148
rect 380124 3136 380130 3188
rect 380894 3136 380900 3188
rect 380952 3176 380958 3188
rect 388438 3176 388444 3188
rect 380952 3148 388444 3176
rect 380952 3136 380958 3148
rect 388438 3136 388444 3148
rect 388496 3136 388502 3188
rect 389818 3136 389824 3188
rect 389876 3176 389882 3188
rect 409598 3176 409604 3188
rect 389876 3148 409604 3176
rect 389876 3136 389882 3148
rect 409598 3136 409604 3148
rect 409656 3136 409662 3188
rect 468478 3136 468484 3188
rect 468536 3176 468542 3188
rect 479334 3176 479340 3188
rect 468536 3148 479340 3176
rect 468536 3136 468542 3148
rect 479334 3136 479340 3148
rect 479392 3136 479398 3188
rect 301958 3068 301964 3120
rect 302016 3108 302022 3120
rect 338298 3108 338304 3120
rect 302016 3080 338304 3108
rect 302016 3068 302022 3080
rect 338298 3068 338304 3080
rect 338356 3068 338362 3120
rect 369854 3068 369860 3120
rect 369912 3108 369918 3120
rect 376570 3108 376576 3120
rect 369912 3080 376576 3108
rect 369912 3068 369918 3080
rect 376570 3068 376576 3080
rect 376628 3068 376634 3120
rect 391842 3108 391848 3120
rect 379486 3080 391848 3108
rect 318518 3000 318524 3052
rect 318576 3040 318582 3052
rect 343818 3040 343824 3052
rect 318576 3012 343824 3040
rect 318576 3000 318582 3012
rect 343818 3000 343824 3012
rect 343876 3000 343882 3052
rect 350442 3000 350448 3052
rect 350500 3040 350506 3052
rect 354674 3040 354680 3052
rect 350500 3012 354680 3040
rect 350500 3000 350506 3012
rect 354674 3000 354680 3012
rect 354732 3000 354738 3052
rect 360378 3000 360384 3052
rect 360436 3040 360442 3052
rect 365806 3040 365812 3052
rect 360436 3012 365812 3040
rect 360436 3000 360442 3012
rect 365806 3000 365812 3012
rect 365864 3000 365870 3052
rect 373258 3000 373264 3052
rect 373316 3040 373322 3052
rect 379486 3040 379514 3080
rect 391842 3068 391848 3080
rect 391900 3068 391906 3120
rect 465718 3068 465724 3120
rect 465776 3108 465782 3120
rect 468662 3108 468668 3120
rect 465776 3080 468668 3108
rect 465776 3068 465782 3080
rect 468662 3068 468668 3080
rect 468720 3068 468726 3120
rect 373316 3012 379514 3040
rect 373316 3000 373322 3012
rect 380158 2932 380164 2984
rect 380216 2972 380222 2984
rect 382366 2972 382372 2984
rect 380216 2944 382372 2972
rect 380216 2932 380222 2944
rect 382366 2932 382372 2944
rect 382424 2932 382430 2984
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 328460 700952 328512 701004
rect 413652 700952 413704 701004
rect 218980 700884 219032 700936
rect 338764 700884 338816 700936
rect 202788 700816 202840 700868
rect 337384 700816 337436 700868
rect 322940 700748 322992 700800
rect 478512 700748 478564 700800
rect 154120 700680 154172 700732
rect 344284 700680 344336 700732
rect 137836 700612 137888 700664
rect 342904 700612 342956 700664
rect 317420 700544 317472 700596
rect 543464 700544 543516 700596
rect 89168 700476 89220 700528
rect 349804 700476 349856 700528
rect 72976 700408 73028 700460
rect 348424 700408 348476 700460
rect 24308 700340 24360 700392
rect 355324 700340 355376 700392
rect 8116 700272 8168 700324
rect 353944 700272 353996 700324
rect 325700 700204 325752 700256
rect 397460 700204 397512 700256
rect 267648 700136 267700 700188
rect 336004 700136 336056 700188
rect 333980 700068 334032 700120
rect 348792 700068 348844 700120
rect 310520 696940 310572 696992
rect 580172 696940 580224 696992
rect 311900 683204 311952 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 361580 683136 361632 683188
rect 309140 670760 309192 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 364432 670692 364484 670744
rect 3424 656888 3476 656940
rect 362960 656888 363012 656940
rect 305000 643084 305052 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 367100 632068 367152 632120
rect 306380 630640 306432 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 369860 618264 369912 618316
rect 303620 616836 303672 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 368480 605820 368532 605872
rect 299572 590656 299624 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 372620 579640 372672 579692
rect 302240 576852 302292 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 375380 565836 375432 565888
rect 298100 563048 298152 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 374000 553392 374052 553444
rect 295340 536800 295392 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 376760 527144 376812 527196
rect 296720 524424 296772 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 380992 514768 381044 514820
rect 293316 510620 293368 510672
rect 580172 510620 580224 510672
rect 276020 502392 276072 502444
rect 579252 502392 579304 502444
rect 270500 502324 270552 502376
rect 579160 502324 579212 502376
rect 330852 502188 330904 502240
rect 364340 502188 364392 502240
rect 299480 502120 299532 502172
rect 335544 502120 335596 502172
rect 325608 502052 325660 502104
rect 429200 502052 429252 502104
rect 234620 501984 234672 502036
rect 340880 501984 340932 502036
rect 322112 501916 322164 501968
rect 462320 501916 462372 501968
rect 320088 501848 320140 501900
rect 494060 501848 494112 501900
rect 169760 501780 169812 501832
rect 346032 501780 346084 501832
rect 315120 501712 315172 501764
rect 558920 501712 558972 501764
rect 104900 501644 104952 501696
rect 351276 501644 351328 501696
rect 40040 501576 40092 501628
rect 356520 501576 356572 501628
rect 265992 501168 266044 501220
rect 579068 501168 579120 501220
rect 260564 501100 260616 501152
rect 578976 501100 579028 501152
rect 255228 501032 255280 501084
rect 578884 501032 578936 501084
rect 3056 500964 3108 501016
rect 358728 500964 358780 501016
rect 336004 500896 336056 500948
rect 337292 500896 337344 500948
rect 337384 500896 337436 500948
rect 342536 500896 342588 500948
rect 348424 500896 348476 500948
rect 353300 500896 353352 500948
rect 355324 500896 355376 500948
rect 360200 500896 360252 500948
rect 338764 500828 338816 500880
rect 344284 500828 344336 500880
rect 353944 500488 353996 500540
rect 358268 500488 358320 500540
rect 342904 500420 342956 500472
rect 347964 500420 348016 500472
rect 349804 500420 349856 500472
rect 354772 500420 354824 500472
rect 282920 500352 282972 500404
rect 339040 500352 339092 500404
rect 344376 500352 344428 500404
rect 349528 500352 349580 500404
rect 358728 500352 358780 500404
rect 379520 500352 379572 500404
rect 234344 500284 234396 500336
rect 409144 500284 409196 500336
rect 316868 500216 316920 500268
rect 527180 500216 527232 500268
rect 267648 500148 267700 500200
rect 578056 500148 578108 500200
rect 3240 500080 3292 500132
rect 382832 500080 382884 500132
rect 4068 500012 4120 500064
rect 384580 500012 384632 500064
rect 3332 499944 3384 499996
rect 386604 499944 386656 499996
rect 3976 499876 4028 499928
rect 388168 499876 388220 499928
rect 3792 499808 3844 499860
rect 389916 499808 389968 499860
rect 3884 499740 3936 499792
rect 391940 499740 391992 499792
rect 3700 499672 3752 499724
rect 393412 499672 393464 499724
rect 3516 499604 3568 499656
rect 395160 499604 395212 499656
rect 3608 499536 3660 499588
rect 396908 499536 396960 499588
rect 233700 499060 233752 499112
rect 402152 499060 402204 499112
rect 234436 498992 234488 499044
rect 405740 498992 405792 499044
rect 234528 498924 234580 498976
rect 407396 498924 407448 498976
rect 234160 498856 234212 498908
rect 411260 498856 411312 498908
rect 234252 498788 234304 498840
rect 412824 498788 412876 498840
rect 288808 498720 288860 498772
rect 580908 498720 580960 498772
rect 274548 498652 274600 498704
rect 577320 498652 577372 498704
rect 272984 498584 273036 498636
rect 577412 498584 577464 498636
rect 269488 498516 269540 498568
rect 578148 498516 578200 498568
rect 264244 498448 264296 498500
rect 577964 498448 578016 498500
rect 258908 498380 258960 498432
rect 577780 498380 577832 498432
rect 250168 498312 250220 498364
rect 574836 498312 574888 498364
rect 253664 498244 253716 498296
rect 577688 498244 577740 498296
rect 248098 498176 248150 498228
rect 577504 498176 577556 498228
rect 278228 497428 278280 497480
rect 279976 497428 280028 497480
rect 281540 497428 281592 497480
rect 283472 497428 283524 497480
rect 285220 497428 285272 497480
rect 286876 497428 286928 497480
rect 290556 497428 290608 497480
rect 292304 497428 292356 497480
rect 580172 497292 580224 497344
rect 580080 497224 580132 497276
rect 580724 497156 580776 497208
rect 580816 497088 580868 497140
rect 580632 497020 580684 497072
rect 580448 496952 580500 497004
rect 580540 496884 580592 496936
rect 580356 496816 580408 496868
rect 235080 338240 235132 338292
rect 235080 337968 235132 338020
rect 314706 337764 314758 337816
rect 314936 337764 314988 337816
rect 259460 336744 259512 336796
rect 259828 336744 259880 336796
rect 307944 336744 307996 336796
rect 308128 336744 308180 336796
rect 321560 336744 321612 336796
rect 321836 336744 321888 336796
rect 173164 336676 173216 336728
rect 270224 336676 270276 336728
rect 274640 336676 274692 336728
rect 275100 336676 275152 336728
rect 305000 336676 305052 336728
rect 339592 336676 339644 336728
rect 354680 336676 354732 336728
rect 354956 336676 355008 336728
rect 360108 336676 360160 336728
rect 360844 336676 360896 336728
rect 369768 336676 369820 336728
rect 373264 336676 373316 336728
rect 373356 336676 373408 336728
rect 378140 336676 378192 336728
rect 378508 336676 378560 336728
rect 380256 336676 380308 336728
rect 386328 336676 386380 336728
rect 411904 336676 411956 336728
rect 414020 336676 414072 336728
rect 414388 336676 414440 336728
rect 426440 336676 426492 336728
rect 427176 336676 427228 336728
rect 428648 336676 428700 336728
rect 451924 336676 451976 336728
rect 163504 336608 163556 336660
rect 267832 336608 267884 336660
rect 298100 336608 298152 336660
rect 337108 336608 337160 336660
rect 360016 336608 360068 336660
rect 362960 336608 363012 336660
rect 373724 336608 373776 336660
rect 400772 336608 400824 336660
rect 433524 336608 433576 336660
rect 458824 336608 458876 336660
rect 153844 336540 153896 336592
rect 265348 336540 265400 336592
rect 291200 336540 291252 336592
rect 328920 336540 328972 336592
rect 149704 336472 149756 336524
rect 264060 336472 264112 336524
rect 287060 336472 287112 336524
rect 333520 336540 333572 336592
rect 345388 336540 345440 336592
rect 353392 336540 353444 336592
rect 364984 336540 365036 336592
rect 377404 336540 377456 336592
rect 388444 336540 388496 336592
rect 416044 336540 416096 336592
rect 434628 336540 434680 336592
rect 472624 336540 472676 336592
rect 145564 336404 145616 336456
rect 261668 336404 261720 336456
rect 284300 336404 284352 336456
rect 332232 336472 332284 336524
rect 366456 336472 366508 336524
rect 379980 336472 380032 336524
rect 389732 336472 389784 336524
rect 433984 336472 434036 336524
rect 331864 336404 331916 336456
rect 345020 336404 345072 336456
rect 375288 336404 375340 336456
rect 402244 336404 402296 336456
rect 426624 336404 426676 336456
rect 475384 336404 475436 336456
rect 45560 336336 45612 336388
rect 250720 336336 250772 336388
rect 262956 336336 263008 336388
rect 315212 336336 315264 336388
rect 316040 336336 316092 336388
rect 343180 336336 343232 336388
rect 368572 336336 368624 336388
rect 384304 336336 384356 336388
rect 394608 336336 394660 336388
rect 460204 336336 460256 336388
rect 38660 336268 38712 336320
rect 248420 336268 248472 336320
rect 264244 336268 264296 336320
rect 318892 336268 318944 336320
rect 328920 336268 328972 336320
rect 334716 336268 334768 336320
rect 31760 336200 31812 336252
rect 245844 336200 245896 336252
rect 273628 336200 273680 336252
rect 328736 336200 328788 336252
rect 24860 336132 24912 336184
rect 243452 336132 243504 336184
rect 261484 336132 261536 336184
rect 319720 336132 319772 336184
rect 327356 336132 327408 336184
rect 347320 336268 347372 336320
rect 369860 336268 369912 336320
rect 388444 336268 388496 336320
rect 393320 336268 393372 336320
rect 460940 336268 460992 336320
rect 334992 336200 335044 336252
rect 347780 336200 347832 336252
rect 371056 336200 371108 336252
rect 396080 336200 396132 336252
rect 399392 336200 399444 336252
rect 468484 336200 468536 336252
rect 334900 336132 334952 336184
rect 346860 336132 346912 336184
rect 372988 336132 373040 336184
rect 393964 336132 394016 336184
rect 395988 336132 396040 336184
rect 465724 336132 465776 336184
rect 15200 336064 15252 336116
rect 240140 336064 240192 336116
rect 269120 336064 269172 336116
rect 327448 336064 327500 336116
rect 334624 336064 334676 336116
rect 349528 336064 349580 336116
rect 377956 336064 378008 336116
rect 405004 336064 405056 336116
rect 416688 336064 416740 336116
rect 528560 336064 528612 336116
rect 5540 335996 5592 336048
rect 236920 335996 236972 336048
rect 266360 335996 266412 336048
rect 326160 335996 326212 336048
rect 331220 335996 331272 336048
rect 348516 335996 348568 336048
rect 366824 335996 366876 336048
rect 374736 335996 374788 336048
rect 376576 335996 376628 336048
rect 406568 335996 406620 336048
rect 418896 335996 418948 336048
rect 535460 335996 535512 336048
rect 177304 335928 177356 335980
rect 271420 335928 271472 335980
rect 307760 335928 307812 335980
rect 340420 335928 340472 335980
rect 373908 335928 373960 335980
rect 181444 335860 181496 335912
rect 273812 335860 273864 335912
rect 311900 335860 311952 335912
rect 342260 335860 342312 335912
rect 370964 335860 371016 335912
rect 374644 335860 374696 335912
rect 380072 335928 380124 335980
rect 406384 335928 406436 335980
rect 426348 335928 426400 335980
rect 447784 335928 447836 335980
rect 398104 335860 398156 335912
rect 412824 335860 412876 335912
rect 434076 335860 434128 335912
rect 188344 335792 188396 335844
rect 276388 335792 276440 335844
rect 318800 335792 318852 335844
rect 344468 335792 344520 335844
rect 362132 335792 362184 335844
rect 363604 335792 363656 335844
rect 376668 335792 376720 335844
rect 391204 335792 391256 335844
rect 421380 335792 421432 335844
rect 440884 335792 440936 335844
rect 236644 335724 236696 335776
rect 277584 335724 277636 335776
rect 326344 335724 326396 335776
rect 338120 335724 338172 335776
rect 375472 335724 375524 335776
rect 389824 335724 389876 335776
rect 431040 335724 431092 335776
rect 450544 335724 450596 335776
rect 260104 335656 260156 335708
rect 294972 335656 295024 335708
rect 325976 335656 326028 335708
rect 334900 335656 334952 335708
rect 374276 335656 374328 335708
rect 387156 335656 387208 335708
rect 423772 335656 423824 335708
rect 440976 335656 441028 335708
rect 329104 335588 329156 335640
rect 339132 335588 339184 335640
rect 333244 335520 333296 335572
rect 334992 335520 335044 335572
rect 371884 335384 371936 335436
rect 376024 335384 376076 335436
rect 353944 335316 353996 335368
rect 356060 335316 356112 335368
rect 266636 330760 266688 330812
rect 266912 330760 266964 330812
rect 291476 330760 291528 330812
rect 292764 330760 292816 330812
rect 301044 330760 301096 330812
rect 320364 330760 320416 330812
rect 291476 330556 291528 330608
rect 292764 330556 292816 330608
rect 301044 330556 301096 330608
rect 320364 330556 320416 330608
rect 234804 330488 234856 330540
rect 235356 330488 235408 330540
rect 238760 330488 238812 330540
rect 239772 330488 239824 330540
rect 240232 330488 240284 330540
rect 240968 330488 241020 330540
rect 244280 330488 244332 330540
rect 244648 330488 244700 330540
rect 245844 330488 245896 330540
rect 246672 330488 246724 330540
rect 249892 330488 249944 330540
rect 250352 330488 250404 330540
rect 252560 330488 252612 330540
rect 253572 330488 253624 330540
rect 255504 330488 255556 330540
rect 256424 330488 256476 330540
rect 256792 330488 256844 330540
rect 257620 330488 257672 330540
rect 258172 330488 258224 330540
rect 258816 330488 258868 330540
rect 259552 330488 259604 330540
rect 260012 330488 260064 330540
rect 262220 330488 262272 330540
rect 262864 330488 262916 330540
rect 267832 330488 267884 330540
rect 268568 330488 268620 330540
rect 270592 330488 270644 330540
rect 271052 330488 271104 330540
rect 271880 330488 271932 330540
rect 272616 330488 272668 330540
rect 273536 330488 273588 330540
rect 274272 330488 274324 330540
rect 276204 330488 276256 330540
rect 276664 330488 276716 330540
rect 278780 330488 278832 330540
rect 279148 330488 279200 330540
rect 280252 330488 280304 330540
rect 280712 330488 280764 330540
rect 283012 330488 283064 330540
rect 283564 330488 283616 330540
rect 284392 330488 284444 330540
rect 284760 330488 284812 330540
rect 285772 330488 285824 330540
rect 286048 330488 286100 330540
rect 287244 330488 287296 330540
rect 287612 330488 287664 330540
rect 288440 330488 288492 330540
rect 288900 330488 288952 330540
rect 289820 330488 289872 330540
rect 290464 330488 290516 330540
rect 291384 330488 291436 330540
rect 292120 330488 292172 330540
rect 292672 330488 292724 330540
rect 293316 330488 293368 330540
rect 294052 330488 294104 330540
rect 294512 330488 294564 330540
rect 296812 330488 296864 330540
rect 297364 330488 297416 330540
rect 298192 330488 298244 330540
rect 298560 330488 298612 330540
rect 299572 330488 299624 330540
rect 300216 330488 300268 330540
rect 300952 330488 301004 330540
rect 301412 330488 301464 330540
rect 311992 330488 312044 330540
rect 312360 330488 312412 330540
rect 313372 330488 313424 330540
rect 314016 330488 314068 330540
rect 314752 330488 314804 330540
rect 315672 330488 315724 330540
rect 316224 330488 316276 330540
rect 316868 330488 316920 330540
rect 317420 330488 317472 330540
rect 318064 330488 318116 330540
rect 320272 330488 320324 330540
rect 320916 330488 320968 330540
rect 321652 330488 321704 330540
rect 322112 330488 322164 330540
rect 324320 330488 324372 330540
rect 325332 330488 325384 330540
rect 327172 330488 327224 330540
rect 327816 330488 327868 330540
rect 328552 330488 328604 330540
rect 329472 330488 329524 330540
rect 340972 330488 341024 330540
rect 341616 330488 341668 330540
rect 345296 330488 345348 330540
rect 346032 330488 346084 330540
rect 349344 330488 349396 330540
rect 349712 330488 349764 330540
rect 360292 330488 360344 330540
rect 360660 330488 360712 330540
rect 363052 330488 363104 330540
rect 363328 330488 363380 330540
rect 367192 330488 367244 330540
rect 367928 330488 367980 330540
rect 379612 330488 379664 330540
rect 380164 330488 380216 330540
rect 382464 330488 382516 330540
rect 383016 330488 383068 330540
rect 383660 330488 383712 330540
rect 384580 330488 384632 330540
rect 386512 330488 386564 330540
rect 387432 330488 387484 330540
rect 410064 330488 410116 330540
rect 410984 330488 411036 330540
rect 411260 330488 411312 330540
rect 411812 330488 411864 330540
rect 414112 330488 414164 330540
rect 414664 330488 414716 330540
rect 427820 330488 427872 330540
rect 428832 330488 428884 330540
rect 429200 330488 429252 330540
rect 430028 330488 430080 330540
rect 430580 330488 430632 330540
rect 431224 330488 431276 330540
rect 234712 330420 234764 330472
rect 235724 330420 235776 330472
rect 244372 330420 244424 330472
rect 245016 330420 245068 330472
rect 255320 330420 255372 330472
rect 255964 330420 256016 330472
rect 259644 330420 259696 330472
rect 260472 330420 260524 330472
rect 262312 330420 262364 330472
rect 263324 330420 263376 330472
rect 276112 330420 276164 330472
rect 277124 330420 277176 330472
rect 280344 330420 280396 330472
rect 281172 330420 281224 330472
rect 284484 330420 284536 330472
rect 285220 330420 285272 330472
rect 287152 330420 287204 330472
rect 288072 330420 288124 330472
rect 288532 330420 288584 330472
rect 289268 330420 289320 330472
rect 298284 330420 298336 330472
rect 299020 330420 299072 330472
rect 312084 330420 312136 330472
rect 312820 330420 312872 330472
rect 317512 330420 317564 330472
rect 318432 330420 318484 330472
rect 360200 330420 360252 330472
rect 361120 330420 361172 330472
rect 379704 330420 379756 330472
rect 380532 330420 380584 330472
rect 382280 330420 382332 330472
rect 383384 330420 383436 330472
rect 409880 330420 409932 330472
rect 410616 330420 410668 330472
rect 411352 330420 411404 330472
rect 412180 330420 412232 330472
rect 414204 330420 414256 330472
rect 415032 330420 415084 330472
rect 430672 330420 430724 330472
rect 431684 330420 431736 330472
rect 349252 330216 349304 330268
rect 350080 330216 350132 330268
rect 258080 330080 258132 330132
rect 258448 330080 258500 330132
rect 299480 330080 299532 330132
rect 299848 330080 299900 330132
rect 253940 329944 253992 329996
rect 254768 329944 254820 329996
rect 295340 329944 295392 329996
rect 296168 329944 296220 329996
rect 416872 329672 416924 329724
rect 417884 329672 417936 329724
rect 387800 329536 387852 329588
rect 388628 329536 388680 329588
rect 256700 329128 256752 329180
rect 257252 329128 257304 329180
rect 313280 328720 313332 328772
rect 313648 328720 313700 328772
rect 365720 328720 365772 328772
rect 366916 328720 366968 328772
rect 283104 328448 283156 328500
rect 284024 328448 284076 328500
rect 363052 328312 363104 328364
rect 363880 328312 363932 328364
rect 289912 327904 289964 327956
rect 290924 327904 290976 327956
rect 329840 327768 329892 327820
rect 330208 327768 330260 327820
rect 260932 327496 260984 327548
rect 261300 327496 261352 327548
rect 408500 327292 408552 327344
rect 409328 327292 409380 327344
rect 296904 327224 296956 327276
rect 297824 327224 297876 327276
rect 325792 326884 325844 326936
rect 326620 326884 326672 326936
rect 285680 326816 285732 326868
rect 286416 326816 286468 326868
rect 329932 326816 329984 326868
rect 330668 326816 330720 326868
rect 419724 326816 419776 326868
rect 280160 326680 280212 326732
rect 280528 326680 280580 326732
rect 309140 326680 309192 326732
rect 309416 326680 309468 326732
rect 419724 326612 419776 326664
rect 396356 326476 396408 326528
rect 396540 326476 396592 326528
rect 303620 326408 303672 326460
rect 304724 326408 304776 326460
rect 305276 326408 305328 326460
rect 305460 326408 305512 326460
rect 306564 326408 306616 326460
rect 307944 326408 307996 326460
rect 308772 326408 308824 326460
rect 310612 326408 310664 326460
rect 311624 326408 311676 326460
rect 335544 326408 335596 326460
rect 335820 326408 335872 326460
rect 352012 326408 352064 326460
rect 352932 326408 352984 326460
rect 397644 326408 397696 326460
rect 398380 326408 398432 326460
rect 404544 326408 404596 326460
rect 405280 326408 405332 326460
rect 303804 326340 303856 326392
rect 304264 326340 304316 326392
rect 305092 326340 305144 326392
rect 305920 326340 305972 326392
rect 307852 326340 307904 326392
rect 308312 326340 308364 326392
rect 309232 326340 309284 326392
rect 309968 326340 310020 326392
rect 310520 326340 310572 326392
rect 311164 326340 311216 326392
rect 332692 326340 332744 326392
rect 333060 326340 333112 326392
rect 335360 326340 335412 326392
rect 335912 326340 335964 326392
rect 338212 326340 338264 326392
rect 338764 326340 338816 326392
rect 350540 326340 350592 326392
rect 351368 326340 351420 326392
rect 351920 326340 351972 326392
rect 352564 326340 352616 326392
rect 353484 326340 353536 326392
rect 354220 326340 354272 326392
rect 354772 326340 354824 326392
rect 355416 326340 355468 326392
rect 389364 326340 389416 326392
rect 390284 326340 390336 326392
rect 394700 326340 394752 326392
rect 395160 326340 395212 326392
rect 396172 326340 396224 326392
rect 396816 326340 396868 326392
rect 397460 326340 397512 326392
rect 398012 326340 398064 326392
rect 398840 326340 398892 326392
rect 399576 326340 399628 326392
rect 400220 326340 400272 326392
rect 401232 326340 401284 326392
rect 402980 326340 403032 326392
rect 403716 326340 403768 326392
rect 404360 326340 404412 326392
rect 404912 326340 404964 326392
rect 405924 326340 405976 326392
rect 406476 326340 406528 326392
rect 407212 326340 407264 326392
rect 408132 326340 408184 326392
rect 418160 326340 418212 326392
rect 419080 326340 419132 326392
rect 419632 326340 419684 326392
rect 420276 326340 420328 326392
rect 420920 326340 420972 326392
rect 421564 326340 421616 326392
rect 422300 326340 422352 326392
rect 423128 326340 423180 326392
rect 242992 326204 243044 326256
rect 243820 326204 243872 326256
rect 306564 326204 306616 326256
rect 335544 326204 335596 326256
rect 336372 326204 336424 326256
rect 400404 326204 400456 326256
rect 400588 326204 400640 326256
rect 401600 325728 401652 325780
rect 402428 325728 402480 325780
rect 577320 325456 577372 325508
rect 580448 325456 580500 325508
rect 390652 325320 390704 325372
rect 391480 325320 391532 325372
rect 400312 324232 400364 324284
rect 400864 324232 400916 324284
rect 306472 323552 306524 323604
rect 306656 323552 306708 323604
rect 352104 323552 352156 323604
rect 352288 323552 352340 323604
rect 422392 323552 422444 323604
rect 422576 323552 422628 323604
rect 425060 323416 425112 323468
rect 425612 323416 425664 323468
rect 390560 323008 390612 323060
rect 391112 323008 391164 323060
rect 306380 322736 306432 322788
rect 307116 322736 307168 322788
rect 389180 322464 389232 322516
rect 389916 322464 389968 322516
rect 423680 322464 423732 322516
rect 424784 322464 424836 322516
rect 423772 322056 423824 322108
rect 424324 322056 424376 322108
rect 403072 321648 403124 321700
rect 403256 321648 403308 321700
rect 419540 319200 419592 319252
rect 419816 319200 419868 319252
rect 3516 306280 3568 306332
rect 233700 306280 233752 306332
rect 577412 299412 577464 299464
rect 579620 299412 579672 299464
rect 3056 293904 3108 293956
rect 233792 293904 233844 293956
rect 578148 273164 578200 273216
rect 579896 273164 579948 273216
rect 3148 255212 3200 255264
rect 234528 255212 234580 255264
rect 578056 245556 578108 245608
rect 579620 245556 579672 245608
rect 3516 241408 3568 241460
rect 234436 241408 234488 241460
rect 577964 233180 578016 233232
rect 579804 233180 579856 233232
rect 3332 215228 3384 215280
rect 234344 215228 234396 215280
rect 577872 206932 577924 206984
rect 579988 206932 580040 206984
rect 3056 202784 3108 202836
rect 234252 202784 234304 202836
rect 577780 193128 577832 193180
rect 579620 193128 579672 193180
rect 3516 188980 3568 189032
rect 234160 188980 234212 189032
rect 3240 164160 3292 164212
rect 234068 164160 234120 164212
rect 577688 153144 577740 153196
rect 580632 153144 580684 153196
rect 3516 150356 3568 150408
rect 235080 150356 235132 150408
rect 3516 137912 3568 137964
rect 233976 137912 234028 137964
rect 577504 112956 577556 113008
rect 580356 112956 580408 113008
rect 3148 111732 3200 111784
rect 233884 111732 233936 111784
rect 574836 100648 574888 100700
rect 580172 100648 580224 100700
rect 577596 73108 577648 73160
rect 579712 73108 579764 73160
rect 574744 60664 574796 60716
rect 580172 60664 580224 60716
rect 74540 20204 74592 20256
rect 259644 20204 259696 20256
rect 70400 20136 70452 20188
rect 259736 20136 259788 20188
rect 67640 20068 67692 20120
rect 258264 20068 258316 20120
rect 63500 20000 63552 20052
rect 256884 20000 256936 20052
rect 60740 19932 60792 19984
rect 255596 19932 255648 19984
rect 187700 19252 187752 19304
rect 299664 19252 299716 19304
rect 151820 19184 151872 19236
rect 287428 19184 287480 19236
rect 121460 19116 121512 19168
rect 276204 19116 276256 19168
rect 118700 19048 118752 19100
rect 274824 19048 274876 19100
rect 114560 18980 114612 19032
rect 273536 18980 273588 19032
rect 56600 18912 56652 18964
rect 254124 18912 254176 18964
rect 52460 18844 52512 18896
rect 252836 18844 252888 18896
rect 49700 18776 49752 18828
rect 251364 18776 251416 18828
rect 44180 18708 44232 18760
rect 249892 18708 249944 18760
rect 41420 18640 41472 18692
rect 248604 18640 248656 18692
rect 37280 18572 37332 18624
rect 247224 18572 247276 18624
rect 191840 18504 191892 18556
rect 301044 18504 301096 18556
rect 194600 18436 194652 18488
rect 301136 18436 301188 18488
rect 198740 18368 198792 18420
rect 302424 18368 302476 18420
rect 208400 17892 208452 17944
rect 306564 17892 306616 17944
rect 204260 17824 204312 17876
rect 305276 17824 305328 17876
rect 201500 17756 201552 17808
rect 303896 17756 303948 17808
rect 197360 17688 197412 17740
rect 302332 17688 302384 17740
rect 153200 17620 153252 17672
rect 287244 17620 287296 17672
rect 150440 17552 150492 17604
rect 285680 17552 285732 17604
rect 151912 17484 151964 17536
rect 287336 17484 287388 17536
rect 149060 17416 149112 17468
rect 285772 17416 285824 17468
rect 146300 17348 146352 17400
rect 284484 17348 284536 17400
rect 147680 17280 147732 17332
rect 285864 17280 285916 17332
rect 143540 17212 143592 17264
rect 284576 17212 284628 17264
rect 211160 17144 211212 17196
rect 308128 17144 308180 17196
rect 224960 17076 225012 17128
rect 312176 17076 312228 17128
rect 227720 17008 227772 17060
rect 313464 17008 313516 17060
rect 164424 16532 164476 16584
rect 291476 16532 291528 16584
rect 161296 16464 161348 16516
rect 290096 16464 290148 16516
rect 143632 16396 143684 16448
rect 283104 16396 283156 16448
rect 125600 16328 125652 16380
rect 277492 16328 277544 16380
rect 123024 16260 123076 16312
rect 276112 16260 276164 16312
rect 119896 16192 119948 16244
rect 276296 16192 276348 16244
rect 116400 16124 116452 16176
rect 274732 16124 274784 16176
rect 112352 16056 112404 16108
rect 273444 16056 273496 16108
rect 34520 15988 34572 16040
rect 245844 15988 245896 16040
rect 30840 15920 30892 15972
rect 245752 15920 245804 15972
rect 27712 15852 27764 15904
rect 244464 15852 244516 15904
rect 168380 15784 168432 15836
rect 292764 15784 292816 15836
rect 171968 15716 172020 15768
rect 294144 15716 294196 15768
rect 221096 15648 221148 15700
rect 310796 15648 310848 15700
rect 98184 15104 98236 15156
rect 267832 15104 267884 15156
rect 93860 15036 93912 15088
rect 266728 15036 266780 15088
rect 91560 14968 91612 15020
rect 266636 14968 266688 15020
rect 87512 14900 87564 14952
rect 265072 14900 265124 14952
rect 84200 14832 84252 14884
rect 263692 14832 263744 14884
rect 80888 14764 80940 14816
rect 262496 14764 262548 14816
rect 77392 14696 77444 14748
rect 260932 14696 260984 14748
rect 73344 14628 73396 14680
rect 259552 14628 259604 14680
rect 69848 14560 69900 14612
rect 258172 14560 258224 14612
rect 66720 14492 66772 14544
rect 256792 14492 256844 14544
rect 63224 14424 63276 14476
rect 255504 14424 255556 14476
rect 102232 14356 102284 14408
rect 269396 14356 269448 14408
rect 105728 14288 105780 14340
rect 270592 14288 270644 14340
rect 109040 14220 109092 14272
rect 272064 14220 272116 14272
rect 108120 13744 108172 13796
rect 271972 13744 272024 13796
rect 404544 13744 404596 13796
rect 497096 13744 497148 13796
rect 104072 13676 104124 13728
rect 270684 13676 270736 13728
rect 405924 13676 405976 13728
rect 500592 13676 500644 13728
rect 100760 13608 100812 13660
rect 269304 13608 269356 13660
rect 407396 13608 407448 13660
rect 503720 13608 503772 13660
rect 97448 13540 97500 13592
rect 267924 13540 267976 13592
rect 408684 13540 408736 13592
rect 507216 13540 507268 13592
rect 93952 13472 94004 13524
rect 266544 13472 266596 13524
rect 410156 13472 410208 13524
rect 511264 13472 511316 13524
rect 59360 13404 59412 13456
rect 255412 13404 255464 13456
rect 411444 13404 411496 13456
rect 514760 13404 514812 13456
rect 56048 13336 56100 13388
rect 254032 13336 254084 13388
rect 414296 13336 414348 13388
rect 521660 13336 521712 13388
rect 52552 13268 52604 13320
rect 252744 13268 252796 13320
rect 414204 13268 414256 13320
rect 525432 13268 525484 13320
rect 48504 13200 48556 13252
rect 251272 13200 251324 13252
rect 417056 13200 417108 13252
rect 532056 13200 532108 13252
rect 44272 13132 44324 13184
rect 249984 13132 250036 13184
rect 422484 13132 422536 13184
rect 546500 13132 546552 13184
rect 40224 13064 40276 13116
rect 248512 13064 248564 13116
rect 429384 13064 429436 13116
rect 567568 13064 567620 13116
rect 110420 12996 110472 13048
rect 273352 12996 273404 13048
rect 403256 12996 403308 13048
rect 493048 12996 493100 13048
rect 156144 12928 156196 12980
rect 288624 12928 288676 12980
rect 390744 12928 390796 12980
rect 454040 12928 454092 12980
rect 160100 12860 160152 12912
rect 290004 12860 290056 12912
rect 219992 12384 220044 12436
rect 310704 12384 310756 12436
rect 397644 12384 397696 12436
rect 476488 12384 476540 12436
rect 216864 12316 216916 12368
rect 309324 12316 309376 12368
rect 400496 12316 400548 12368
rect 481732 12316 481784 12368
rect 213368 12248 213420 12300
rect 308036 12248 308088 12300
rect 403164 12248 403216 12300
rect 489920 12248 489972 12300
rect 209780 12180 209832 12232
rect 306472 12180 306524 12232
rect 404452 12180 404504 12232
rect 494704 12180 494756 12232
rect 206192 12112 206244 12164
rect 305184 12112 305236 12164
rect 202696 12044 202748 12096
rect 303804 12044 303856 12096
rect 145472 11976 145524 12028
rect 284392 11976 284444 12028
rect 316224 12112 316276 12164
rect 418252 12112 418304 12164
rect 534448 12112 534500 12164
rect 419724 12044 419776 12096
rect 538220 12044 538272 12096
rect 421012 11976 421064 12028
rect 541992 11976 542044 12028
rect 142160 11908 142212 11960
rect 283012 11908 283064 11960
rect 316132 11908 316184 11960
rect 421104 11908 421156 11960
rect 545488 11908 545540 11960
rect 138848 11840 138900 11892
rect 281724 11840 281776 11892
rect 422392 11840 422444 11892
rect 547880 11840 547932 11892
rect 135260 11772 135312 11824
rect 280344 11772 280396 11824
rect 423864 11772 423916 11824
rect 551008 11772 551060 11824
rect 131304 11704 131356 11756
rect 280436 11704 280488 11756
rect 425152 11704 425204 11756
rect 554780 11704 554832 11756
rect 143540 11636 143592 11688
rect 144736 11636 144788 11688
rect 223580 11636 223632 11688
rect 310612 11636 310664 11688
rect 396448 11636 396500 11688
rect 473452 11636 473504 11688
rect 226340 11568 226392 11620
rect 312084 11568 312136 11620
rect 396356 11568 396408 11620
rect 469864 11568 469916 11620
rect 231032 11500 231084 11552
rect 313372 11500 313424 11552
rect 394792 11500 394844 11552
rect 465632 11500 465684 11552
rect 173900 10956 173952 11008
rect 294052 10956 294104 11008
rect 393412 10956 393464 11008
rect 463976 10956 464028 11008
rect 170312 10888 170364 10940
rect 292672 10888 292724 10940
rect 394700 10888 394752 10940
rect 467472 10888 467524 10940
rect 167184 10820 167236 10872
rect 291384 10820 291436 10872
rect 396264 10820 396316 10872
rect 470600 10820 470652 10872
rect 163412 10752 163464 10804
rect 289912 10752 289964 10804
rect 397552 10752 397604 10804
rect 474096 10752 474148 10804
rect 158904 10684 158956 10736
rect 288532 10684 288584 10736
rect 398932 10684 398984 10736
rect 478144 10684 478196 10736
rect 155408 10616 155460 10668
rect 287152 10616 287204 10668
rect 400404 10616 400456 10668
rect 482376 10616 482428 10668
rect 89904 10548 89956 10600
rect 265164 10548 265216 10600
rect 398840 10548 398892 10600
rect 480536 10548 480588 10600
rect 86408 10480 86460 10532
rect 263784 10480 263836 10532
rect 400312 10480 400364 10532
rect 484032 10480 484084 10532
rect 83280 10412 83332 10464
rect 262312 10412 262364 10464
rect 401692 10412 401744 10464
rect 486424 10412 486476 10464
rect 79232 10344 79284 10396
rect 262404 10344 262456 10396
rect 401784 10344 401836 10396
rect 487160 10344 487212 10396
rect 75920 10276 75972 10328
rect 261024 10276 261076 10328
rect 403072 10276 403124 10328
rect 490656 10276 490708 10328
rect 176660 10208 176712 10260
rect 295524 10208 295576 10260
rect 392124 10208 392176 10260
rect 459928 10208 459980 10260
rect 180984 10140 181036 10192
rect 297088 10140 297140 10192
rect 390652 10140 390704 10192
rect 456892 10140 456944 10192
rect 184940 10072 184992 10124
rect 298376 10072 298428 10124
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 222752 9596 222804 9648
rect 310520 9596 310572 9648
rect 387892 9596 387944 9648
rect 446220 9596 446272 9648
rect 219256 9528 219308 9580
rect 309232 9528 309284 9580
rect 316040 9528 316092 9580
rect 316316 9528 316368 9580
rect 389272 9528 389324 9580
rect 449808 9528 449860 9580
rect 215668 9460 215720 9512
rect 307944 9460 307996 9512
rect 315948 9460 316000 9512
rect 316224 9460 316276 9512
rect 389364 9460 389416 9512
rect 453304 9460 453356 9512
rect 137652 9392 137704 9444
rect 281632 9392 281684 9444
rect 422300 9392 422352 9444
rect 549076 9392 549128 9444
rect 37188 9324 37240 9376
rect 247132 9324 247184 9376
rect 277124 9324 277176 9376
rect 330024 9324 330076 9376
rect 423772 9324 423824 9376
rect 552664 9324 552716 9376
rect 33600 9256 33652 9308
rect 245936 9256 245988 9308
rect 262956 9256 263008 9308
rect 324596 9256 324648 9308
rect 425060 9256 425112 9308
rect 556160 9256 556212 9308
rect 30104 9188 30156 9240
rect 244372 9188 244424 9240
rect 259460 9188 259512 9240
rect 323124 9188 323176 9240
rect 426532 9188 426584 9240
rect 559748 9188 559800 9240
rect 26516 9120 26568 9172
rect 242992 9120 243044 9172
rect 255872 9120 255924 9172
rect 321836 9120 321888 9172
rect 428004 9120 428056 9172
rect 563244 9120 563296 9172
rect 21824 9052 21876 9104
rect 241704 9052 241756 9104
rect 252376 9052 252428 9104
rect 321744 9052 321796 9104
rect 429292 9052 429344 9104
rect 566832 9052 566884 9104
rect 8760 8984 8812 9036
rect 237472 8984 237524 9036
rect 242072 8984 242124 9036
rect 317696 8984 317748 9036
rect 430764 8984 430816 9036
rect 570328 8984 570380 9036
rect 4068 8916 4120 8968
rect 236092 8916 236144 8968
rect 238116 8916 238168 8968
rect 316408 8916 316460 8968
rect 430672 8916 430724 8968
rect 573916 8916 573968 8968
rect 226432 8848 226484 8900
rect 311992 8848 312044 8900
rect 386696 8848 386748 8900
rect 442632 8848 442684 8900
rect 229836 8780 229888 8832
rect 313280 8780 313332 8832
rect 385132 8780 385184 8832
rect 439136 8780 439188 8832
rect 233424 8712 233476 8764
rect 314844 8712 314896 8764
rect 383844 8712 383896 8764
rect 435548 8712 435600 8764
rect 183744 8236 183796 8288
rect 296904 8236 296956 8288
rect 404360 8236 404412 8288
rect 495900 8236 495952 8288
rect 180248 8168 180300 8220
rect 296996 8168 297048 8220
rect 405832 8168 405884 8220
rect 499396 8168 499448 8220
rect 176752 8100 176804 8152
rect 295432 8100 295484 8152
rect 407304 8100 407356 8152
rect 502984 8100 503036 8152
rect 173072 8032 173124 8084
rect 294236 8032 294288 8084
rect 408592 8032 408644 8084
rect 506480 8032 506532 8084
rect 169576 7964 169628 8016
rect 292580 7964 292632 8016
rect 409972 7964 410024 8016
rect 510068 7964 510120 8016
rect 162492 7896 162544 7948
rect 289820 7896 289872 7948
rect 290740 7896 290792 7948
rect 320364 7896 320416 7948
rect 410064 7896 410116 7948
rect 513564 7896 513616 7948
rect 157800 7828 157852 7880
rect 288440 7828 288492 7880
rect 288532 7828 288584 7880
rect 328552 7828 328604 7880
rect 411352 7828 411404 7880
rect 517152 7828 517204 7880
rect 130568 7760 130620 7812
rect 278964 7760 279016 7812
rect 286600 7760 286652 7812
rect 332692 7760 332744 7812
rect 412732 7760 412784 7812
rect 520740 7760 520792 7812
rect 126980 7692 127032 7744
rect 277584 7692 277636 7744
rect 283104 7692 283156 7744
rect 331496 7692 331548 7744
rect 414112 7692 414164 7744
rect 524236 7692 524288 7744
rect 128176 7624 128228 7676
rect 278872 7624 278924 7676
rect 279516 7624 279568 7676
rect 329932 7624 329984 7676
rect 415492 7624 415544 7676
rect 527824 7624 527876 7676
rect 69112 7556 69164 7608
rect 258080 7556 258132 7608
rect 272432 7556 272484 7608
rect 328644 7556 328696 7608
rect 416964 7556 417016 7608
rect 531320 7556 531372 7608
rect 187332 7488 187384 7540
rect 298284 7488 298336 7540
rect 402980 7488 403032 7540
rect 492312 7488 492364 7540
rect 190828 7420 190880 7472
rect 299572 7420 299624 7472
rect 401600 7420 401652 7472
rect 488816 7420 488868 7472
rect 194416 7352 194468 7404
rect 300952 7352 301004 7404
rect 400220 7352 400272 7404
rect 485228 7352 485280 7404
rect 62028 6808 62080 6860
rect 255320 6808 255372 6860
rect 271236 6808 271288 6860
rect 327172 6808 327224 6860
rect 387800 6808 387852 6860
rect 448612 6808 448664 6860
rect 58440 6740 58492 6792
rect 253940 6740 253992 6792
rect 268844 6740 268896 6792
rect 327264 6740 327316 6792
rect 389180 6740 389232 6792
rect 452108 6740 452160 6792
rect 54944 6672 54996 6724
rect 252560 6672 252612 6724
rect 265348 6672 265400 6724
rect 325884 6672 325936 6724
rect 390560 6672 390612 6724
rect 455696 6672 455748 6724
rect 51356 6604 51408 6656
rect 252652 6604 252704 6656
rect 261760 6604 261812 6656
rect 324504 6604 324556 6656
rect 392032 6604 392084 6656
rect 459192 6604 459244 6656
rect 47860 6536 47912 6588
rect 251180 6536 251232 6588
rect 258264 6536 258316 6588
rect 323032 6536 323084 6588
rect 393320 6536 393372 6588
rect 462780 6536 462832 6588
rect 17040 6468 17092 6520
rect 240324 6468 240376 6520
rect 254676 6468 254728 6520
rect 321652 6468 321704 6520
rect 383752 6468 383804 6520
rect 12348 6400 12400 6452
rect 238944 6400 238996 6452
rect 251180 6400 251232 6452
rect 320272 6400 320324 6452
rect 433984 6468 434036 6520
rect 434076 6468 434128 6520
rect 518348 6468 518400 6520
rect 7656 6332 7708 6384
rect 237380 6332 237432 6384
rect 239312 6332 239364 6384
rect 316132 6332 316184 6384
rect 379704 6332 379756 6384
rect 424968 6332 425020 6384
rect 427912 6332 427964 6384
rect 562048 6400 562100 6452
rect 436744 6332 436796 6384
rect 565636 6332 565688 6384
rect 2872 6264 2924 6316
rect 234712 6264 234764 6316
rect 240508 6264 240560 6316
rect 317604 6264 317656 6316
rect 380992 6264 381044 6316
rect 427268 6264 427320 6316
rect 429200 6264 429252 6316
rect 569132 6264 569184 6316
rect 1676 6196 1728 6248
rect 234804 6196 234856 6248
rect 235816 6196 235868 6248
rect 314752 6196 314804 6248
rect 381084 6196 381136 6248
rect 428464 6196 428516 6248
rect 430580 6196 430632 6248
rect 572720 6196 572772 6248
rect 572 6128 624 6180
rect 234620 6128 234672 6180
rect 237012 6128 237064 6180
rect 316040 6128 316092 6180
rect 432052 6128 432104 6180
rect 576308 6128 576360 6180
rect 65524 6060 65576 6112
rect 256700 6060 256752 6112
rect 285404 6060 285456 6112
rect 332784 6060 332836 6112
rect 386512 6060 386564 6112
rect 445024 6060 445076 6112
rect 136456 5992 136508 6044
rect 281540 5992 281592 6044
rect 288992 5992 289044 6044
rect 334072 5992 334124 6044
rect 386604 5992 386656 6044
rect 441528 5992 441580 6044
rect 140044 5924 140096 5976
rect 282920 5924 282972 5976
rect 309876 5924 309928 5976
rect 334164 5924 334216 5976
rect 385040 5924 385092 5976
rect 437940 5924 437992 5976
rect 234620 5856 234672 5908
rect 262864 5856 262916 5908
rect 382556 5856 382608 5908
rect 430856 5856 430908 5908
rect 382464 5788 382516 5840
rect 432052 5788 432104 5840
rect 427820 5720 427872 5772
rect 436744 5720 436796 5772
rect 210976 5448 211028 5500
rect 306380 5448 306432 5500
rect 407212 5448 407264 5500
rect 505376 5448 505428 5500
rect 85672 5380 85724 5432
rect 149704 5380 149756 5432
rect 207388 5380 207440 5432
rect 305092 5380 305144 5432
rect 324412 5380 324464 5432
rect 345296 5380 345348 5432
rect 408500 5380 408552 5432
rect 508872 5380 508924 5432
rect 89168 5312 89220 5364
rect 153844 5312 153896 5364
rect 203892 5312 203944 5364
rect 303620 5312 303672 5364
rect 317328 5312 317380 5364
rect 343732 5312 343784 5364
rect 409880 5312 409932 5364
rect 512460 5312 512512 5364
rect 78588 5244 78640 5296
rect 145564 5244 145616 5296
rect 196808 5244 196860 5296
rect 302240 5244 302292 5296
rect 313832 5244 313884 5296
rect 342352 5244 342404 5296
rect 411260 5244 411312 5296
rect 515956 5244 516008 5296
rect 96252 5176 96304 5228
rect 163504 5176 163556 5228
rect 193220 5176 193272 5228
rect 300860 5176 300912 5228
rect 310244 5176 310296 5228
rect 341064 5176 341116 5228
rect 367284 5176 367336 5228
rect 387156 5176 387208 5228
rect 412640 5176 412692 5228
rect 519544 5176 519596 5228
rect 121092 5108 121144 5160
rect 188344 5108 188396 5160
rect 189724 5108 189776 5160
rect 299480 5108 299532 5160
rect 306748 5108 306800 5160
rect 339592 5108 339644 5160
rect 371332 5108 371384 5160
rect 400128 5108 400180 5160
rect 414020 5108 414072 5160
rect 523040 5108 523092 5160
rect 114008 5040 114060 5092
rect 181444 5040 181496 5092
rect 186136 5040 186188 5092
rect 298192 5040 298244 5092
rect 303160 5040 303212 5092
rect 338212 5040 338264 5092
rect 367100 5040 367152 5092
rect 367284 5040 367336 5092
rect 374000 5040 374052 5092
rect 407212 5040 407264 5092
rect 415400 5040 415452 5092
rect 526628 5040 526680 5092
rect 103336 4972 103388 5024
rect 173164 4972 173216 5024
rect 182548 4972 182600 5024
rect 296812 4972 296864 5024
rect 299664 4972 299716 5024
rect 336924 4972 336976 5024
rect 375380 4972 375432 5024
rect 410800 4972 410852 5024
rect 416780 4972 416832 5024
rect 530124 4972 530176 5024
rect 106924 4904 106976 4956
rect 177304 4904 177356 4956
rect 179052 4904 179104 4956
rect 295340 4904 295392 4956
rect 296076 4904 296128 4956
rect 335544 4904 335596 4956
rect 376760 4904 376812 4956
rect 414296 4904 414348 4956
rect 418160 4904 418212 4956
rect 537208 4904 537260 4956
rect 132960 4836 133012 4888
rect 280160 4836 280212 4888
rect 292580 4836 292632 4888
rect 335636 4836 335688 4888
rect 378232 4836 378284 4888
rect 417884 4836 417936 4888
rect 419632 4836 419684 4888
rect 540796 4836 540848 4888
rect 129372 4768 129424 4820
rect 278780 4768 278832 4820
rect 281908 4768 281960 4820
rect 331404 4768 331456 4820
rect 378324 4768 378376 4820
rect 420184 4768 420236 4820
rect 420920 4768 420972 4820
rect 544384 4768 544436 4820
rect 214472 4700 214524 4752
rect 307852 4700 307904 4752
rect 407120 4700 407172 4752
rect 501788 4700 501840 4752
rect 218060 4632 218112 4684
rect 309140 4632 309192 4684
rect 405740 4632 405792 4684
rect 498200 4632 498252 4684
rect 175464 4564 175516 4616
rect 260104 4564 260156 4616
rect 299296 4564 299348 4616
rect 329840 4564 329892 4616
rect 379612 4564 379664 4616
rect 423772 4564 423824 4616
rect 298008 4496 298060 4548
rect 324320 4496 324372 4548
rect 379520 4496 379572 4548
rect 421380 4496 421432 4548
rect 299388 4428 299440 4480
rect 324228 4428 324280 4480
rect 378140 4428 378192 4480
rect 418988 4428 419040 4480
rect 301504 4360 301556 4412
rect 325792 4360 325844 4412
rect 328736 4292 328788 4344
rect 176660 4156 176712 4208
rect 177856 4156 177908 4208
rect 226340 4156 226392 4208
rect 227536 4156 227588 4208
rect 99840 4088 99892 4140
rect 269212 4088 269264 4140
rect 274824 4088 274876 4140
rect 311440 4088 311492 4140
rect 340880 4088 340932 4140
rect 342168 4088 342220 4140
rect 352104 4088 352156 4140
rect 363236 4088 363288 4140
rect 367100 4088 367152 4140
rect 367192 4088 367244 4140
rect 378784 4088 378836 4140
rect 92756 4020 92808 4072
rect 266452 4020 266504 4072
rect 267740 4020 267792 4072
rect 301504 4020 301556 4072
rect 309048 4020 309100 4072
rect 340788 4020 340840 4072
rect 340972 4020 341024 4072
rect 82084 3952 82136 4004
rect 262220 3952 262272 4004
rect 264152 3952 264204 4004
rect 299388 3952 299440 4004
rect 317880 3952 317932 4004
rect 322940 3952 322992 4004
rect 338672 3952 338724 4004
rect 350724 3952 350776 4004
rect 351644 4020 351696 4072
rect 354772 4020 354824 4072
rect 360844 4020 360896 4072
rect 364616 4020 364668 4072
rect 365720 4020 365772 4072
rect 400864 4156 400916 4208
rect 383660 4088 383712 4140
rect 384764 4020 384816 4072
rect 388352 4088 388404 4140
rect 402520 4088 402572 4140
rect 403624 4088 403676 4140
rect 405004 4088 405056 4140
rect 411904 4088 411956 4140
rect 411996 4088 412048 4140
rect 440332 4088 440384 4140
rect 440976 4088 441028 4140
rect 550272 4088 550324 4140
rect 352196 3952 352248 4004
rect 360292 3952 360344 4004
rect 367008 3952 367060 4004
rect 368480 3952 368532 4004
rect 43076 3884 43128 3936
rect 248696 3884 248748 3936
rect 276020 3884 276072 3936
rect 288532 3884 288584 3936
rect 294880 3884 294932 3936
rect 335360 3884 335412 3936
rect 336280 3884 336332 3936
rect 349252 3884 349304 3936
rect 363144 3884 363196 3936
rect 377404 3952 377456 4004
rect 378876 3952 378928 4004
rect 378968 3952 379020 4004
rect 388260 3952 388312 4004
rect 391204 4020 391256 4072
rect 413100 4020 413152 4072
rect 416044 4020 416096 4072
rect 447416 4020 447468 4072
rect 447784 4020 447836 4072
rect 557356 4020 557408 4072
rect 393136 3952 393188 4004
rect 402704 3952 402756 4004
rect 404820 3952 404872 4004
rect 405740 3952 405792 4004
rect 472256 3952 472308 4004
rect 472624 3952 472676 4004
rect 582196 3952 582248 4004
rect 35992 3816 36044 3868
rect 247040 3816 247092 3868
rect 248788 3816 248840 3868
rect 290740 3816 290792 3868
rect 293684 3816 293736 3868
rect 335452 3816 335504 3868
rect 337476 3816 337528 3868
rect 350632 3816 350684 3868
rect 363052 3816 363104 3868
rect 370872 3816 370924 3868
rect 374092 3816 374144 3868
rect 382280 3884 382332 3936
rect 433248 3884 433300 3936
rect 433892 3884 433944 3936
rect 450912 3884 450964 3936
rect 451924 3884 451976 3936
rect 564440 3884 564492 3936
rect 390652 3816 390704 3868
rect 391940 3816 391992 3868
rect 458088 3816 458140 3868
rect 458824 3816 458876 3868
rect 578608 3816 578660 3868
rect 28908 3748 28960 3800
rect 244280 3748 244332 3800
rect 245200 3748 245252 3800
rect 264244 3748 264296 3800
rect 280712 3748 280764 3800
rect 331312 3748 331364 3800
rect 332692 3748 332744 3800
rect 349528 3748 349580 3800
rect 363328 3748 363380 3800
rect 363696 3748 363748 3800
rect 367100 3748 367152 3800
rect 375288 3748 375340 3800
rect 376024 3748 376076 3800
rect 398932 3748 398984 3800
rect 402612 3748 402664 3800
rect 408408 3748 408460 3800
rect 409144 3748 409196 3800
rect 415492 3748 415544 3800
rect 419540 3748 419592 3800
rect 539600 3748 539652 3800
rect 24216 3680 24268 3732
rect 243084 3680 243136 3732
rect 257068 3680 257120 3732
rect 317880 3680 317932 3732
rect 20628 3612 20680 3664
rect 241612 3612 241664 3664
rect 253480 3612 253532 3664
rect 321560 3680 321612 3732
rect 330392 3680 330444 3732
rect 347872 3680 347924 3732
rect 360200 3680 360252 3732
rect 19432 3544 19484 3596
rect 241520 3544 241572 3596
rect 249984 3544 250036 3596
rect 320180 3612 320232 3664
rect 325608 3612 325660 3664
rect 346492 3612 346544 3664
rect 349252 3612 349304 3664
rect 354864 3612 354916 3664
rect 361580 3612 361632 3664
rect 365812 3680 365864 3732
rect 381176 3680 381228 3732
rect 388444 3680 388496 3732
rect 393044 3680 393096 3732
rect 393136 3680 393188 3732
rect 436744 3680 436796 3732
rect 450544 3680 450596 3732
rect 571524 3680 571576 3732
rect 318892 3544 318944 3596
rect 323308 3544 323360 3596
rect 345204 3544 345256 3596
rect 368204 3612 368256 3664
rect 370872 3612 370924 3664
rect 376484 3612 376536 3664
rect 376576 3612 376628 3664
rect 394240 3612 394292 3664
rect 394332 3612 394384 3664
rect 401324 3612 401376 3664
rect 406384 3612 406436 3664
rect 369400 3544 369452 3596
rect 371240 3544 371292 3596
rect 397736 3544 397788 3596
rect 398104 3544 398156 3596
rect 402704 3544 402756 3596
rect 406476 3544 406528 3596
rect 411904 3544 411956 3596
rect 412088 3612 412140 3664
rect 416688 3612 416740 3664
rect 423680 3612 423732 3664
rect 553768 3612 553820 3664
rect 422576 3544 422628 3596
rect 426440 3544 426492 3596
rect 560852 3544 560904 3596
rect 14740 3476 14792 3528
rect 238760 3476 238812 3528
rect 246396 3476 246448 3528
rect 322112 3476 322164 3528
rect 345112 3476 345164 3528
rect 11152 3408 11204 3460
rect 238852 3408 238904 3460
rect 242900 3408 242952 3460
rect 317420 3408 317472 3460
rect 329196 3408 329248 3460
rect 333244 3408 333296 3460
rect 333888 3408 333940 3460
rect 334624 3408 334676 3460
rect 344560 3408 344612 3460
rect 352012 3476 352064 3528
rect 352840 3476 352892 3528
rect 353944 3476 353996 3528
rect 355232 3476 355284 3528
rect 356244 3476 356296 3528
rect 357532 3476 357584 3528
rect 358728 3476 358780 3528
rect 358912 3476 358964 3528
rect 361120 3476 361172 3528
rect 364340 3476 364392 3528
rect 377680 3476 377732 3528
rect 380256 3476 380308 3528
rect 388352 3476 388404 3528
rect 388444 3476 388496 3528
rect 426164 3476 426216 3528
rect 431960 3476 432012 3528
rect 575112 3476 575164 3528
rect 44180 3340 44232 3392
rect 45100 3340 45152 3392
rect 52460 3340 52512 3392
rect 53380 3340 53432 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 110512 3272 110564 3324
rect 271880 3340 271932 3392
rect 278320 3340 278372 3392
rect 299296 3340 299348 3392
rect 315028 3340 315080 3392
rect 342444 3340 342496 3392
rect 117596 3272 117648 3324
rect 274640 3272 274692 3324
rect 300768 3272 300820 3324
rect 326436 3272 326488 3324
rect 335084 3272 335136 3324
rect 349344 3408 349396 3460
rect 364432 3408 364484 3460
rect 348056 3340 348108 3392
rect 353484 3340 353536 3392
rect 361672 3340 361724 3392
rect 371700 3340 371752 3392
rect 382372 3408 382424 3460
rect 429660 3408 429712 3460
rect 433340 3408 433392 3460
rect 581000 3408 581052 3460
rect 379980 3340 380032 3392
rect 380072 3340 380124 3392
rect 395344 3340 395396 3392
rect 396172 3340 396224 3392
rect 405740 3340 405792 3392
rect 440884 3340 440936 3392
rect 543188 3340 543240 3392
rect 346952 3272 347004 3324
rect 353392 3272 353444 3324
rect 354036 3272 354088 3324
rect 356152 3272 356204 3324
rect 367284 3272 367336 3324
rect 385960 3272 386012 3324
rect 387064 3272 387116 3324
rect 124680 3204 124732 3256
rect 236644 3204 236696 3256
rect 260656 3204 260708 3256
rect 298008 3204 298060 3256
rect 304356 3204 304408 3256
rect 329104 3204 329156 3256
rect 339868 3204 339920 3256
rect 350540 3204 350592 3256
rect 363696 3204 363748 3256
rect 372896 3204 372948 3256
rect 374736 3204 374788 3256
rect 383568 3204 383620 3256
rect 384304 3204 384356 3256
rect 389456 3204 389508 3256
rect 397460 3272 397512 3324
rect 475752 3272 475804 3324
rect 406016 3204 406068 3256
rect 460204 3204 460256 3256
rect 465172 3204 465224 3256
rect 475384 3204 475436 3256
rect 558552 3272 558604 3324
rect 247592 3136 247644 3188
rect 261484 3136 261536 3188
rect 290188 3136 290240 3188
rect 309876 3136 309928 3188
rect 320916 3136 320968 3188
rect 331864 3136 331916 3188
rect 343364 3136 343416 3188
rect 351920 3136 351972 3188
rect 359004 3136 359056 3188
rect 362316 3136 362368 3188
rect 363604 3136 363656 3188
rect 370596 3136 370648 3188
rect 374644 3136 374696 3188
rect 380072 3136 380124 3188
rect 380900 3136 380952 3188
rect 388444 3136 388496 3188
rect 389824 3136 389876 3188
rect 409604 3136 409656 3188
rect 468484 3136 468536 3188
rect 479340 3136 479392 3188
rect 301964 3068 302016 3120
rect 338304 3068 338356 3120
rect 369860 3068 369912 3120
rect 376576 3068 376628 3120
rect 318524 3000 318576 3052
rect 343824 3000 343876 3052
rect 350448 3000 350500 3052
rect 354680 3000 354732 3052
rect 360384 3000 360436 3052
rect 365812 3000 365864 3052
rect 373264 3000 373316 3052
rect 391848 3068 391900 3120
rect 465724 3068 465776 3120
rect 468668 3068 468720 3120
rect 380164 2932 380216 2984
rect 382372 2932 382424 2984
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 40052 501634 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 104912 501702 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 137848 700670 137876 703520
rect 154132 700738 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 169772 501838 169800 702406
rect 202800 700874 202828 703520
rect 218992 700942 219020 703520
rect 218980 700936 219032 700942
rect 218980 700878 219032 700884
rect 202788 700868 202840 700874
rect 202788 700810 202840 700816
rect 234632 502042 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700194 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 700188 267700 700194
rect 267648 700130 267700 700136
rect 276020 502444 276072 502450
rect 276020 502386 276072 502392
rect 270500 502376 270552 502382
rect 270500 502318 270552 502324
rect 234620 502036 234672 502042
rect 234620 501978 234672 501984
rect 169760 501832 169812 501838
rect 169760 501774 169812 501780
rect 104900 501696 104952 501702
rect 104900 501638 104952 501644
rect 40040 501628 40092 501634
rect 40040 501570 40092 501576
rect 265992 501220 266044 501226
rect 265992 501162 266044 501168
rect 260564 501152 260616 501158
rect 260564 501094 260616 501100
rect 255228 501084 255280 501090
rect 255228 501026 255280 501032
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 500440 3478 500449
rect 3422 500375 3478 500384
rect 3240 500132 3292 500138
rect 3240 500074 3292 500080
rect 3252 475697 3280 500074
rect 3332 499996 3384 500002
rect 3332 499938 3384 499944
rect 3238 475688 3294 475697
rect 3238 475623 3294 475632
rect 3344 462641 3372 499938
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 6497 3464 500375
rect 234344 500336 234396 500342
rect 234344 500278 234396 500284
rect 4068 500064 4120 500070
rect 4068 500006 4120 500012
rect 3976 499928 4028 499934
rect 3976 499870 4028 499876
rect 3792 499860 3844 499866
rect 3792 499802 3844 499808
rect 3700 499724 3752 499730
rect 3700 499666 3752 499672
rect 3516 499656 3568 499662
rect 3516 499598 3568 499604
rect 3528 345409 3556 499598
rect 3608 499588 3660 499594
rect 3608 499530 3660 499536
rect 3620 358465 3648 499530
rect 3712 371385 3740 499666
rect 3804 397497 3832 499802
rect 3884 499792 3936 499798
rect 3884 499734 3936 499740
rect 3896 410553 3924 499734
rect 3988 423609 4016 499870
rect 4080 449585 4108 500006
rect 233700 499112 233752 499118
rect 233700 499054 233752 499060
rect 4066 449576 4122 449585
rect 4066 449511 4122 449520
rect 3974 423600 4030 423609
rect 3974 423535 4030 423544
rect 3882 410544 3938 410553
rect 3882 410479 3938 410488
rect 3790 397488 3846 397497
rect 3790 397423 3846 397432
rect 3698 371376 3754 371385
rect 3698 371311 3754 371320
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 173164 336728 173216 336734
rect 173164 336670 173216 336676
rect 163504 336660 163556 336666
rect 163504 336602 163556 336608
rect 153844 336592 153896 336598
rect 153844 336534 153896 336540
rect 149704 336524 149756 336530
rect 149704 336466 149756 336472
rect 145564 336456 145616 336462
rect 145564 336398 145616 336404
rect 45560 336388 45612 336394
rect 45560 336330 45612 336336
rect 38660 336320 38712 336326
rect 38660 336262 38712 336268
rect 31760 336252 31812 336258
rect 31760 336194 31812 336200
rect 24860 336184 24912 336190
rect 24860 336126 24912 336132
rect 15200 336116 15252 336122
rect 15200 336058 15252 336064
rect 5540 336048 5592 336054
rect 5540 335990 5592 335996
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 5552 16574 5580 335990
rect 9678 18592 9734 18601
rect 9678 18527 9734 18536
rect 5552 16546 6040 16574
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 572 6180 624 6186
rect 572 6122 624 6128
rect 584 480 612 6122
rect 1688 480 1716 6190
rect 2884 480 2912 6258
rect 4080 480 4108 8910
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7668 480 7696 6326
rect 8772 480 8800 8978
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 18527
rect 15212 16574 15240 336058
rect 24872 16574 24900 336126
rect 31772 16574 31800 336194
rect 37280 18624 37332 18630
rect 37280 18566 37332 18572
rect 37292 16574 37320 18566
rect 38672 16574 38700 336262
rect 44180 18760 44232 18766
rect 44180 18702 44232 18708
rect 41420 18692 41472 18698
rect 41420 18634 41472 18640
rect 41432 16574 41460 18634
rect 15212 16546 15976 16574
rect 24872 16546 25360 16574
rect 31772 16546 31984 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 41432 16546 41920 16574
rect 13542 11656 13598 11665
rect 13542 11591 13598 11600
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 12360 480 12388 6394
rect 13556 480 13584 11591
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 480 14780 3470
rect 15948 480 15976 16546
rect 22558 14512 22614 14521
rect 22558 14447 22614 14456
rect 17958 13016 18014 13025
rect 17958 12951 18014 12960
rect 17040 6520 17092 6526
rect 17040 6462 17092 6468
rect 17052 480 17080 6462
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 12951
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19444 480 19472 3538
rect 20640 480 20668 3606
rect 21836 480 21864 9046
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 14447
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24228 480 24256 3674
rect 25332 480 25360 16546
rect 30840 15972 30892 15978
rect 30840 15914 30892 15920
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 26516 9172 26568 9178
rect 26516 9114 26568 9120
rect 26528 480 26556 9114
rect 27724 480 27752 15846
rect 30104 9240 30156 9246
rect 30104 9182 30156 9188
rect 28908 3800 28960 3806
rect 28908 3742 28960 3748
rect 28920 480 28948 3742
rect 30116 480 30144 9182
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 15914
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 34520 16040 34572 16046
rect 34520 15982 34572 15988
rect 33600 9308 33652 9314
rect 33600 9250 33652 9256
rect 33612 480 33640 9250
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 15982
rect 37188 9376 37240 9382
rect 37188 9318 37240 9324
rect 35992 3868 36044 3874
rect 35992 3810 36044 3816
rect 36004 480 36032 3810
rect 37200 480 37228 9318
rect 38396 480 38424 16546
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 40224 13116 40276 13122
rect 40224 13058 40276 13064
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 13058
rect 41892 480 41920 16546
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 43088 480 43116 3878
rect 44192 3398 44220 18702
rect 45572 16574 45600 336330
rect 74540 20256 74592 20262
rect 74540 20198 74592 20204
rect 70400 20188 70452 20194
rect 70400 20130 70452 20136
rect 67640 20120 67692 20126
rect 67640 20062 67692 20068
rect 63500 20052 63552 20058
rect 63500 19994 63552 20000
rect 60740 19984 60792 19990
rect 60740 19926 60792 19932
rect 56600 18964 56652 18970
rect 56600 18906 56652 18912
rect 52460 18896 52512 18902
rect 52460 18838 52512 18844
rect 49700 18828 49752 18834
rect 49700 18770 49752 18776
rect 49712 16574 49740 18770
rect 45572 16546 46704 16574
rect 49712 16546 50200 16574
rect 44272 13184 44324 13190
rect 44272 13126 44324 13132
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44284 480 44312 13126
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45112 354 45140 3334
rect 46676 480 46704 16546
rect 48504 13252 48556 13258
rect 48504 13194 48556 13200
rect 47860 6588 47912 6594
rect 47860 6530 47912 6536
rect 47872 480 47900 6530
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 13194
rect 50172 480 50200 16546
rect 51356 6656 51408 6662
rect 51356 6598 51408 6604
rect 51368 480 51396 6598
rect 52472 3398 52500 18838
rect 56612 16574 56640 18906
rect 60752 16574 60780 19926
rect 63512 16574 63540 19994
rect 56612 16546 56824 16574
rect 60752 16546 60872 16574
rect 63512 16546 64368 16574
rect 56048 13388 56100 13394
rect 56048 13330 56100 13336
rect 52552 13320 52604 13326
rect 52552 13262 52604 13268
rect 52460 3392 52512 3398
rect 52460 3334 52512 3340
rect 52564 480 52592 13262
rect 54944 6724 54996 6730
rect 54944 6666 54996 6672
rect 53380 3392 53432 3398
rect 53380 3334 53432 3340
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3334
rect 54956 480 54984 6666
rect 56060 480 56088 13330
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 59360 13456 59412 13462
rect 59360 13398 59412 13404
rect 58440 6792 58492 6798
rect 58440 6734 58492 6740
rect 58452 480 58480 6734
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 13398
rect 60844 480 60872 16546
rect 63224 14476 63276 14482
rect 63224 14418 63276 14424
rect 62028 6860 62080 6866
rect 62028 6802 62080 6808
rect 62040 480 62068 6802
rect 63236 480 63264 14418
rect 64340 480 64368 16546
rect 66720 14544 66772 14550
rect 66720 14486 66772 14492
rect 65524 6112 65576 6118
rect 65524 6054 65576 6060
rect 65536 480 65564 6054
rect 66732 480 66760 14486
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 20062
rect 70412 16574 70440 20130
rect 74552 16574 74580 20198
rect 121460 19168 121512 19174
rect 121460 19110 121512 19116
rect 118700 19100 118752 19106
rect 118700 19042 118752 19048
rect 114560 19032 114612 19038
rect 114560 18974 114612 18980
rect 114572 16574 114600 18974
rect 118712 16574 118740 19042
rect 121472 16574 121500 19110
rect 143540 17264 143592 17270
rect 140778 17232 140834 17241
rect 143540 17206 143592 17212
rect 140778 17167 140834 17176
rect 140792 16574 140820 17167
rect 70412 16546 71544 16574
rect 74552 16546 75040 16574
rect 114572 16546 114784 16574
rect 118712 16546 118832 16574
rect 121472 16546 122328 16574
rect 140792 16546 141280 16574
rect 69848 14612 69900 14618
rect 69848 14554 69900 14560
rect 69112 7608 69164 7614
rect 69112 7550 69164 7556
rect 69124 480 69152 7550
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 14554
rect 71516 480 71544 16546
rect 73344 14680 73396 14686
rect 73344 14622 73396 14628
rect 72606 10296 72662 10305
rect 72606 10231 72662 10240
rect 72620 480 72648 10231
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 14622
rect 75012 480 75040 16546
rect 112352 16108 112404 16114
rect 112352 16050 112404 16056
rect 98184 15156 98236 15162
rect 98184 15098 98236 15104
rect 93860 15088 93912 15094
rect 93860 15030 93912 15036
rect 91560 15020 91612 15026
rect 91560 14962 91612 14968
rect 87512 14952 87564 14958
rect 87512 14894 87564 14900
rect 84200 14884 84252 14890
rect 84200 14826 84252 14832
rect 80888 14816 80940 14822
rect 80888 14758 80940 14764
rect 77392 14748 77444 14754
rect 77392 14690 77444 14696
rect 75920 10328 75972 10334
rect 75920 10270 75972 10276
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 10270
rect 77404 480 77432 14690
rect 79232 10396 79284 10402
rect 79232 10338 79284 10344
rect 78588 5296 78640 5302
rect 78588 5238 78640 5244
rect 78600 480 78628 5238
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 10338
rect 80900 480 80928 14758
rect 83280 10464 83332 10470
rect 83280 10406 83332 10412
rect 82084 4004 82136 4010
rect 82084 3946 82136 3952
rect 82096 480 82124 3946
rect 83292 480 83320 10406
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 14826
rect 86408 10532 86460 10538
rect 86408 10474 86460 10480
rect 85672 5432 85724 5438
rect 85672 5374 85724 5380
rect 85684 480 85712 5374
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 10474
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 14894
rect 89904 10600 89956 10606
rect 89904 10542 89956 10548
rect 89168 5364 89220 5370
rect 89168 5306 89220 5312
rect 89180 480 89208 5306
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 10542
rect 91572 480 91600 14962
rect 92756 4072 92808 4078
rect 92756 4014 92808 4020
rect 92768 480 92796 4014
rect 93872 3398 93900 15030
rect 97448 13592 97500 13598
rect 97448 13534 97500 13540
rect 93952 13524 94004 13530
rect 93952 13466 94004 13472
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 13466
rect 96252 5228 96304 5234
rect 96252 5170 96304 5176
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 96264 480 96292 5170
rect 97460 480 97488 13534
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 15098
rect 102232 14408 102284 14414
rect 102232 14350 102284 14356
rect 100760 13660 100812 13666
rect 100760 13602 100812 13608
rect 99840 4140 99892 4146
rect 99840 4082 99892 4088
rect 99852 480 99880 4082
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 13602
rect 102244 480 102272 14350
rect 105728 14340 105780 14346
rect 105728 14282 105780 14288
rect 104072 13728 104124 13734
rect 104072 13670 104124 13676
rect 103336 5024 103388 5030
rect 103336 4966 103388 4972
rect 103348 480 103376 4966
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 13670
rect 105740 480 105768 14282
rect 109040 14272 109092 14278
rect 109040 14214 109092 14220
rect 108120 13796 108172 13802
rect 108120 13738 108172 13744
rect 106924 4956 106976 4962
rect 106924 4898 106976 4904
rect 106936 480 106964 4898
rect 108132 480 108160 13738
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 14214
rect 110420 13048 110472 13054
rect 110420 12990 110472 12996
rect 110432 3398 110460 12990
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 110512 3324 110564 3330
rect 110512 3266 110564 3272
rect 110524 480 110552 3266
rect 111628 480 111656 3334
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16050
rect 114008 5092 114060 5098
rect 114008 5034 114060 5040
rect 114020 480 114048 5034
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116400 16176 116452 16182
rect 116400 16118 116452 16124
rect 116412 480 116440 16118
rect 117596 3324 117648 3330
rect 117596 3266 117648 3272
rect 117608 480 117636 3266
rect 118804 480 118832 16546
rect 119896 16244 119948 16250
rect 119896 16186 119948 16192
rect 119908 480 119936 16186
rect 121092 5160 121144 5166
rect 121092 5102 121144 5108
rect 121104 480 121132 5102
rect 122300 480 122328 16546
rect 125600 16380 125652 16386
rect 125600 16322 125652 16328
rect 123024 16312 123076 16318
rect 123024 16254 123076 16260
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16254
rect 124680 3256 124732 3262
rect 124680 3198 124732 3204
rect 124692 480 124720 3198
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 16322
rect 138848 11892 138900 11898
rect 138848 11834 138900 11840
rect 135260 11824 135312 11830
rect 135260 11766 135312 11772
rect 131304 11756 131356 11762
rect 131304 11698 131356 11704
rect 130568 7812 130620 7818
rect 130568 7754 130620 7760
rect 126980 7744 127032 7750
rect 126980 7686 127032 7692
rect 126992 480 127020 7686
rect 128176 7676 128228 7682
rect 128176 7618 128228 7624
rect 128188 480 128216 7618
rect 129372 4820 129424 4826
rect 129372 4762 129424 4768
rect 129384 480 129412 4762
rect 130580 480 130608 7754
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 11698
rect 134154 8936 134210 8945
rect 134154 8871 134210 8880
rect 132960 4888 133012 4894
rect 132960 4830 133012 4836
rect 132972 480 133000 4830
rect 134168 480 134196 8871
rect 135272 480 135300 11766
rect 137652 9444 137704 9450
rect 137652 9386 137704 9392
rect 136456 6044 136508 6050
rect 136456 5986 136508 5992
rect 136468 480 136496 5986
rect 137664 480 137692 9386
rect 138860 480 138888 11834
rect 140044 5976 140096 5982
rect 140044 5918 140096 5924
rect 140056 480 140084 5918
rect 141252 480 141280 16546
rect 142160 11960 142212 11966
rect 142160 11902 142212 11908
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142172 354 142200 11902
rect 143552 11694 143580 17206
rect 143632 16448 143684 16454
rect 143632 16390 143684 16396
rect 143540 11688 143592 11694
rect 143540 11630 143592 11636
rect 143644 6914 143672 16390
rect 145472 12028 145524 12034
rect 145472 11970 145524 11976
rect 144736 11688 144788 11694
rect 144736 11630 144788 11636
rect 143552 6886 143672 6914
rect 143552 480 143580 6886
rect 144748 480 144776 11630
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 11970
rect 145576 5302 145604 336398
rect 149060 17468 149112 17474
rect 149060 17410 149112 17416
rect 146300 17400 146352 17406
rect 146300 17342 146352 17348
rect 146312 16574 146340 17342
rect 147680 17332 147732 17338
rect 147680 17274 147732 17280
rect 147692 16574 147720 17274
rect 149072 16574 149100 17410
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 145564 5296 145616 5302
rect 145564 5238 145616 5244
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 149716 5438 149744 336466
rect 151820 19236 151872 19242
rect 151820 19178 151872 19184
rect 150440 17604 150492 17610
rect 150440 17546 150492 17552
rect 150452 16574 150480 17546
rect 150452 16546 150664 16574
rect 149704 5432 149756 5438
rect 149704 5374 149756 5380
rect 150636 480 150664 16546
rect 151832 9674 151860 19178
rect 153200 17672 153252 17678
rect 153200 17614 153252 17620
rect 151912 17536 151964 17542
rect 151912 17478 151964 17484
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 17478
rect 153212 16574 153240 17614
rect 153212 16546 153792 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 153856 5370 153884 336534
rect 161296 16516 161348 16522
rect 161296 16458 161348 16464
rect 156144 12980 156196 12986
rect 156144 12922 156196 12928
rect 155408 10668 155460 10674
rect 155408 10610 155460 10616
rect 153844 5364 153896 5370
rect 153844 5306 153896 5312
rect 155420 480 155448 10610
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 12922
rect 160100 12912 160152 12918
rect 160100 12854 160152 12860
rect 158904 10736 158956 10742
rect 158904 10678 158956 10684
rect 157800 7880 157852 7886
rect 157800 7822 157852 7828
rect 157812 480 157840 7822
rect 158916 480 158944 10678
rect 160112 480 160140 12854
rect 161308 480 161336 16458
rect 163412 10804 163464 10810
rect 163412 10746 163464 10752
rect 162492 7948 162544 7954
rect 162492 7890 162544 7896
rect 162504 480 162532 7890
rect 163424 3482 163452 10746
rect 163516 5234 163544 336602
rect 164424 16584 164476 16590
rect 164424 16526 164476 16532
rect 163504 5228 163556 5234
rect 163504 5170 163556 5176
rect 163424 3454 163728 3482
rect 163700 480 163728 3454
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 16526
rect 168380 15836 168432 15842
rect 168380 15778 168432 15784
rect 167184 10872 167236 10878
rect 167184 10814 167236 10820
rect 166078 7576 166134 7585
rect 166078 7511 166134 7520
rect 166092 480 166120 7511
rect 167196 480 167224 10814
rect 168392 480 168420 15778
rect 171968 15768 172020 15774
rect 171968 15710 172020 15716
rect 170312 10940 170364 10946
rect 170312 10882 170364 10888
rect 169576 8016 169628 8022
rect 169576 7958 169628 7964
rect 169588 480 169616 7958
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 10882
rect 171980 480 172008 15710
rect 173072 8084 173124 8090
rect 173072 8026 173124 8032
rect 173084 3482 173112 8026
rect 173176 5030 173204 336670
rect 177304 335980 177356 335986
rect 177304 335922 177356 335928
rect 173900 11008 173952 11014
rect 173900 10950 173952 10956
rect 173164 5024 173216 5030
rect 173164 4966 173216 4972
rect 173084 3454 173204 3482
rect 173176 480 173204 3454
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 10950
rect 176660 10260 176712 10266
rect 176660 10202 176712 10208
rect 175464 4616 175516 4622
rect 175464 4558 175516 4564
rect 175476 480 175504 4558
rect 176672 4214 176700 10202
rect 176752 8152 176804 8158
rect 176752 8094 176804 8100
rect 176660 4208 176712 4214
rect 176660 4150 176712 4156
rect 176764 3482 176792 8094
rect 177316 4962 177344 335922
rect 181444 335912 181496 335918
rect 181444 335854 181496 335860
rect 180984 10192 181036 10198
rect 180984 10134 181036 10140
rect 180248 8220 180300 8226
rect 180248 8162 180300 8168
rect 177304 4956 177356 4962
rect 177304 4898 177356 4904
rect 179052 4956 179104 4962
rect 179052 4898 179104 4904
rect 177856 4208 177908 4214
rect 177856 4150 177908 4156
rect 176672 3454 176792 3482
rect 176672 480 176700 3454
rect 177868 480 177896 4150
rect 179064 480 179092 4898
rect 180260 480 180288 8162
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 10134
rect 181456 5098 181484 335854
rect 188344 335844 188396 335850
rect 188344 335786 188396 335792
rect 187700 19304 187752 19310
rect 187700 19246 187752 19252
rect 187712 16574 187740 19246
rect 187712 16546 188292 16574
rect 184940 10124 184992 10130
rect 184940 10066 184992 10072
rect 183744 8288 183796 8294
rect 183744 8230 183796 8236
rect 181444 5092 181496 5098
rect 181444 5034 181496 5040
rect 182548 5024 182600 5030
rect 182548 4966 182600 4972
rect 182560 480 182588 4966
rect 183756 480 183784 8230
rect 184952 480 184980 10066
rect 187332 7540 187384 7546
rect 187332 7482 187384 7488
rect 186136 5092 186188 5098
rect 186136 5034 186188 5040
rect 186148 480 186176 5034
rect 187344 480 187372 7482
rect 188264 3482 188292 16546
rect 188356 5166 188384 335786
rect 233712 306338 233740 499054
rect 234160 498908 234212 498914
rect 234160 498850 234212 498856
rect 233974 498808 234030 498817
rect 233974 498743 234030 498752
rect 233882 497312 233938 497321
rect 233882 497247 233938 497256
rect 233790 496224 233846 496233
rect 233790 496159 233846 496168
rect 233700 306332 233752 306338
rect 233700 306274 233752 306280
rect 233804 293962 233832 496159
rect 233792 293956 233844 293962
rect 233792 293898 233844 293904
rect 233896 111790 233924 497247
rect 233988 137970 234016 498743
rect 234066 497584 234122 497593
rect 234066 497519 234122 497528
rect 234080 164218 234108 497519
rect 234172 189038 234200 498850
rect 234252 498840 234304 498846
rect 234252 498782 234304 498788
rect 234264 202842 234292 498782
rect 234356 215286 234384 500278
rect 235906 500032 235962 500041
rect 235906 499967 235962 499976
rect 234436 499044 234488 499050
rect 234436 498986 234488 498992
rect 234448 241466 234476 498986
rect 234528 498976 234580 498982
rect 234528 498918 234580 498924
rect 234540 255270 234568 498918
rect 235920 498250 235948 499967
rect 246670 499896 246726 499905
rect 246670 499831 246726 499840
rect 241242 499760 241298 499769
rect 241242 499695 241298 499704
rect 235874 498222 235948 498250
rect 239356 498264 239412 498273
rect 235874 497964 235902 498222
rect 239356 498199 239412 498208
rect 239370 497964 239398 498199
rect 241256 497978 241284 499695
rect 244922 498536 244978 498545
rect 244922 498471 244978 498480
rect 242806 498400 242862 498409
rect 242806 498335 242862 498344
rect 241132 497950 241284 497978
rect 242820 497978 242848 498335
rect 244936 497978 244964 498471
rect 246684 497978 246712 499831
rect 250168 498364 250220 498370
rect 250168 498306 250220 498312
rect 248098 498228 248150 498234
rect 248098 498170 248150 498176
rect 242820 497950 242880 497978
rect 244628 497950 244964 497978
rect 246376 497950 246712 497978
rect 248110 497964 248138 498170
rect 250180 497978 250208 498306
rect 253664 498296 253716 498302
rect 253664 498238 253716 498244
rect 253676 497978 253704 498238
rect 255240 497978 255268 501026
rect 258908 498432 258960 498438
rect 258908 498374 258960 498380
rect 258920 497978 258948 498374
rect 260576 497978 260604 501094
rect 264244 498500 264296 498506
rect 264244 498442 264296 498448
rect 264256 497978 264284 498442
rect 266004 497978 266032 501162
rect 267648 500200 267700 500206
rect 267648 500142 267700 500148
rect 267660 497978 267688 500142
rect 269488 498568 269540 498574
rect 269488 498510 269540 498516
rect 269500 497978 269528 498510
rect 249872 497950 250208 497978
rect 253368 497950 253704 497978
rect 255116 497950 255268 497978
rect 258612 497950 258948 497978
rect 260360 497950 260604 497978
rect 263948 497950 264284 497978
rect 265696 497950 266032 497978
rect 267444 497950 267688 497978
rect 269192 497950 269528 497978
rect 270512 497978 270540 502318
rect 274548 498704 274600 498710
rect 274548 498646 274600 498652
rect 272984 498636 273036 498642
rect 272984 498578 273036 498584
rect 272996 497978 273024 498578
rect 274560 497978 274588 498646
rect 270512 497950 270940 497978
rect 272688 497950 273024 497978
rect 274436 497950 274588 497978
rect 276032 497978 276060 502386
rect 282932 500410 282960 702406
rect 298100 563100 298152 563106
rect 298100 563042 298152 563048
rect 295340 536852 295392 536858
rect 295340 536794 295392 536800
rect 293316 510672 293368 510678
rect 293316 510614 293368 510620
rect 282920 500404 282972 500410
rect 282920 500346 282972 500352
rect 288808 498772 288860 498778
rect 288808 498714 288860 498720
rect 288820 497978 288848 498714
rect 276032 497950 276184 497978
rect 288512 497950 288848 497978
rect 293328 497978 293356 510614
rect 295352 497978 295380 536794
rect 296720 524476 296772 524482
rect 296720 524418 296772 524424
rect 296732 518894 296760 524418
rect 298112 518894 298140 563042
rect 296732 518866 296852 518894
rect 298112 518866 298600 518894
rect 296824 497978 296852 518866
rect 298572 497978 298600 518866
rect 299492 502178 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 328460 701004 328512 701010
rect 328460 700946 328512 700952
rect 322940 700800 322992 700806
rect 322940 700742 322992 700748
rect 317420 700596 317472 700602
rect 317420 700538 317472 700544
rect 310520 696992 310572 696998
rect 310520 696934 310572 696940
rect 309140 670812 309192 670818
rect 309140 670754 309192 670760
rect 305000 643136 305052 643142
rect 305000 643078 305052 643084
rect 303620 616888 303672 616894
rect 303620 616830 303672 616836
rect 299572 590708 299624 590714
rect 299572 590650 299624 590656
rect 299584 518894 299612 590650
rect 302240 576904 302292 576910
rect 302240 576846 302292 576852
rect 299584 518866 300348 518894
rect 299480 502172 299532 502178
rect 299480 502114 299532 502120
rect 300320 497978 300348 518866
rect 302252 497978 302280 576846
rect 303632 518894 303660 616830
rect 305012 518894 305040 643078
rect 306380 630692 306432 630698
rect 306380 630634 306432 630640
rect 306392 518894 306420 630634
rect 303632 518866 303844 518894
rect 305012 518866 305592 518894
rect 306392 518866 307340 518894
rect 303816 497978 303844 518866
rect 305564 497978 305592 518866
rect 307312 497978 307340 518866
rect 309152 497978 309180 670754
rect 310532 518894 310560 696934
rect 311900 683256 311952 683262
rect 311900 683198 311952 683204
rect 311912 518894 311940 683198
rect 317432 518894 317460 700538
rect 322952 518894 322980 700742
rect 325700 700256 325752 700262
rect 325700 700198 325752 700204
rect 325712 518894 325740 700198
rect 310532 518866 310928 518894
rect 311912 518866 312676 518894
rect 317432 518866 317920 518894
rect 322952 518866 323164 518894
rect 325712 518866 326660 518894
rect 310900 497978 310928 518866
rect 312648 497978 312676 518866
rect 315120 501764 315172 501770
rect 315120 501706 315172 501712
rect 315132 497978 315160 501706
rect 316868 500268 316920 500274
rect 316868 500210 316920 500216
rect 316880 497978 316908 500210
rect 293328 497950 293756 497978
rect 295352 497950 295504 497978
rect 296824 497950 297252 497978
rect 298572 497950 299000 497978
rect 300320 497950 300748 497978
rect 302252 497950 302496 497978
rect 303816 497950 304244 497978
rect 305564 497950 305992 497978
rect 307312 497950 307740 497978
rect 309152 497950 309488 497978
rect 310900 497950 311328 497978
rect 312648 497950 313076 497978
rect 314824 497950 315160 497978
rect 316572 497950 316908 497978
rect 317892 497978 317920 518866
rect 322112 501968 322164 501974
rect 322112 501910 322164 501916
rect 320088 501900 320140 501906
rect 320088 501842 320140 501848
rect 320100 498250 320128 501842
rect 320054 498222 320128 498250
rect 317892 497950 318320 497978
rect 320054 497964 320082 498222
rect 322124 497978 322152 501910
rect 321816 497950 322152 497978
rect 323136 497978 323164 518866
rect 325608 502104 325660 502110
rect 325608 502046 325660 502052
rect 325620 497978 325648 502046
rect 323136 497950 323564 497978
rect 325312 497950 325648 497978
rect 326632 497978 326660 518866
rect 328472 497978 328500 700946
rect 331232 518894 331260 702986
rect 338764 700936 338816 700942
rect 338764 700878 338816 700884
rect 337384 700868 337436 700874
rect 337384 700810 337436 700816
rect 336004 700188 336056 700194
rect 336004 700130 336056 700136
rect 333980 700120 334032 700126
rect 333980 700062 334032 700068
rect 331232 518866 331904 518894
rect 330852 502240 330904 502246
rect 330852 502182 330904 502188
rect 330864 497978 330892 502182
rect 326632 497950 327060 497978
rect 328472 497950 328808 497978
rect 330556 497950 330892 497978
rect 331876 497978 331904 518866
rect 333992 497978 334020 700062
rect 335544 502172 335596 502178
rect 335544 502114 335596 502120
rect 335556 497978 335584 502114
rect 336016 500954 336044 700130
rect 337396 500954 337424 700810
rect 336004 500948 336056 500954
rect 336004 500890 336056 500896
rect 337292 500948 337344 500954
rect 337292 500890 337344 500896
rect 337384 500948 337436 500954
rect 337384 500890 337436 500896
rect 337304 497978 337332 500890
rect 338776 500886 338804 700878
rect 344284 700732 344336 700738
rect 344284 700674 344336 700680
rect 342904 700664 342956 700670
rect 342904 700606 342956 700612
rect 340880 502036 340932 502042
rect 340880 501978 340932 501984
rect 338764 500880 338816 500886
rect 338764 500822 338816 500828
rect 339040 500404 339092 500410
rect 339040 500346 339092 500352
rect 339052 497978 339080 500346
rect 340892 497978 340920 501978
rect 342536 500948 342588 500954
rect 342536 500890 342588 500896
rect 342548 497978 342576 500890
rect 342916 500478 342944 700606
rect 344296 518894 344324 700674
rect 348424 700460 348476 700466
rect 348424 700402 348476 700408
rect 344296 518866 344416 518894
rect 344284 500880 344336 500886
rect 344284 500822 344336 500828
rect 342904 500472 342956 500478
rect 342904 500414 342956 500420
rect 344296 497978 344324 500822
rect 344388 500410 344416 518866
rect 346032 501832 346084 501838
rect 346032 501774 346084 501780
rect 344376 500404 344428 500410
rect 344376 500346 344428 500352
rect 346044 497978 346072 501774
rect 348436 500954 348464 700402
rect 348804 700126 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 349804 700528 349856 700534
rect 349804 700470 349856 700476
rect 348792 700120 348844 700126
rect 348792 700062 348844 700068
rect 348424 500948 348476 500954
rect 348424 500890 348476 500896
rect 349816 500478 349844 700470
rect 355324 700392 355376 700398
rect 355324 700334 355376 700340
rect 353944 700324 353996 700330
rect 353944 700266 353996 700272
rect 351276 501696 351328 501702
rect 351276 501638 351328 501644
rect 347964 500472 348016 500478
rect 347964 500414 348016 500420
rect 349804 500472 349856 500478
rect 349804 500414 349856 500420
rect 347976 497978 348004 500414
rect 349528 500404 349580 500410
rect 349528 500346 349580 500352
rect 349540 497978 349568 500346
rect 351288 497978 351316 501638
rect 353300 500948 353352 500954
rect 353300 500890 353352 500896
rect 353312 497978 353340 500890
rect 353956 500546 353984 700266
rect 355336 500954 355364 700334
rect 361580 683188 361632 683194
rect 361580 683130 361632 683136
rect 361592 518894 361620 683130
rect 362960 656940 363012 656946
rect 362960 656882 363012 656888
rect 362972 518894 363000 656882
rect 361592 518866 361804 518894
rect 362972 518866 363552 518894
rect 356520 501628 356572 501634
rect 356520 501570 356572 501576
rect 355324 500948 355376 500954
rect 355324 500890 355376 500896
rect 353944 500540 353996 500546
rect 353944 500482 353996 500488
rect 354772 500472 354824 500478
rect 354772 500414 354824 500420
rect 354784 497978 354812 500414
rect 356532 497978 356560 501570
rect 358728 501016 358780 501022
rect 358728 500958 358780 500964
rect 358268 500540 358320 500546
rect 358268 500482 358320 500488
rect 358280 497978 358308 500482
rect 358740 500410 358768 500958
rect 360200 500948 360252 500954
rect 360200 500890 360252 500896
rect 358728 500404 358780 500410
rect 358728 500346 358780 500352
rect 360212 497978 360240 500890
rect 361776 497978 361804 518866
rect 363524 497978 363552 518866
rect 364352 502246 364380 702406
rect 397472 700262 397500 703520
rect 413664 701010 413692 703520
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 364432 670744 364484 670750
rect 364432 670686 364484 670692
rect 364444 518894 364472 670686
rect 367100 632120 367152 632126
rect 367100 632062 367152 632068
rect 364444 518866 365300 518894
rect 364340 502240 364392 502246
rect 364340 502182 364392 502188
rect 365272 497978 365300 518866
rect 367112 497978 367140 632062
rect 369860 618316 369912 618322
rect 369860 618258 369912 618264
rect 368480 605872 368532 605878
rect 368480 605814 368532 605820
rect 368492 518894 368520 605814
rect 369872 518894 369900 618258
rect 372620 579692 372672 579698
rect 372620 579634 372672 579640
rect 368492 518866 368796 518894
rect 369872 518866 370544 518894
rect 368768 497978 368796 518866
rect 370516 497978 370544 518866
rect 372632 497978 372660 579634
rect 375380 565888 375432 565894
rect 375380 565830 375432 565836
rect 374000 553444 374052 553450
rect 374000 553386 374052 553392
rect 374012 497978 374040 553386
rect 375392 518894 375420 565830
rect 376760 527196 376812 527202
rect 376760 527138 376812 527144
rect 376772 518894 376800 527138
rect 375392 518866 375788 518894
rect 376772 518866 377536 518894
rect 375760 497978 375788 518866
rect 377508 497978 377536 518866
rect 380992 514820 381044 514826
rect 380992 514762 381044 514768
rect 379520 500404 379572 500410
rect 379520 500346 379572 500352
rect 379532 497978 379560 500346
rect 381004 497978 381032 514762
rect 429212 502110 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 502104 429252 502110
rect 429200 502046 429252 502052
rect 462332 501974 462360 703520
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 462320 501968 462372 501974
rect 462320 501910 462372 501916
rect 494072 501906 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 501900 494112 501906
rect 494060 501842 494112 501848
rect 431958 500440 432014 500449
rect 431958 500375 432014 500384
rect 409144 500336 409196 500342
rect 398838 500304 398894 500313
rect 409144 500278 409196 500284
rect 398838 500239 398894 500248
rect 382832 500132 382884 500138
rect 382832 500074 382884 500080
rect 382844 497978 382872 500074
rect 384580 500064 384632 500070
rect 384580 500006 384632 500012
rect 384592 497978 384620 500006
rect 386604 499996 386656 500002
rect 386604 499938 386656 499944
rect 386616 497978 386644 499938
rect 388168 499928 388220 499934
rect 388168 499870 388220 499876
rect 388180 497978 388208 499870
rect 389916 499860 389968 499866
rect 389916 499802 389968 499808
rect 389928 497978 389956 499802
rect 391940 499792 391992 499798
rect 391940 499734 391992 499740
rect 391952 497978 391980 499734
rect 393412 499724 393464 499730
rect 393412 499666 393464 499672
rect 393424 497978 393452 499666
rect 395160 499656 395212 499662
rect 395160 499598 395212 499604
rect 395172 497978 395200 499598
rect 396908 499588 396960 499594
rect 396908 499530 396960 499536
rect 396920 497978 396948 499530
rect 398852 497978 398880 500239
rect 403898 500168 403954 500177
rect 403898 500103 403954 500112
rect 402152 499112 402204 499118
rect 402152 499054 402204 499060
rect 402164 497978 402192 499054
rect 403912 497978 403940 500103
rect 405740 499044 405792 499050
rect 405740 498986 405792 498992
rect 405752 497978 405780 498986
rect 407396 498976 407448 498982
rect 407396 498918 407448 498924
rect 407408 497978 407436 498918
rect 409156 497978 409184 500278
rect 411260 498908 411312 498914
rect 411260 498850 411312 498856
rect 411272 497978 411300 498850
rect 412824 498840 412876 498846
rect 412824 498782 412876 498788
rect 416226 498808 416282 498817
rect 412836 497978 412864 498782
rect 416226 498743 416282 498752
rect 416240 497978 416268 498743
rect 421470 498672 421526 498681
rect 421470 498607 421526 498616
rect 421484 497978 421512 498607
rect 431972 497978 432000 500375
rect 527192 500274 527220 703520
rect 543476 700602 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700596 543516 700602
rect 543464 700538 543516 700544
rect 558932 501770 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 579252 502444 579304 502450
rect 579252 502386 579304 502392
rect 579160 502376 579212 502382
rect 579160 502318 579212 502324
rect 558920 501764 558972 501770
rect 558920 501706 558972 501712
rect 579068 501220 579120 501226
rect 579068 501162 579120 501168
rect 578976 501152 579028 501158
rect 578976 501094 579028 501100
rect 578884 501084 578936 501090
rect 578884 501026 578936 501032
rect 527180 500268 527232 500274
rect 527180 500210 527232 500216
rect 578056 500200 578108 500206
rect 578056 500142 578108 500148
rect 436742 500032 436798 500041
rect 436742 499967 436798 499976
rect 331876 497950 332304 497978
rect 333992 497950 334052 497978
rect 335556 497950 335892 497978
rect 337304 497950 337640 497978
rect 339052 497950 339388 497978
rect 340892 497950 341136 497978
rect 342548 497950 342884 497978
rect 344296 497950 344632 497978
rect 346044 497950 346380 497978
rect 347976 497950 348128 497978
rect 349540 497950 349876 497978
rect 351288 497950 351624 497978
rect 353312 497950 353372 497978
rect 354784 497950 355120 497978
rect 356532 497950 356868 497978
rect 358280 497950 358616 497978
rect 360212 497950 360364 497978
rect 361776 497950 362204 497978
rect 363524 497950 363952 497978
rect 365272 497950 365700 497978
rect 367112 497950 367448 497978
rect 368768 497950 369196 497978
rect 370516 497950 370944 497978
rect 372632 497950 372692 497978
rect 374012 497950 374440 497978
rect 375760 497950 376188 497978
rect 377508 497950 377936 497978
rect 379532 497950 379684 497978
rect 381004 497950 381432 497978
rect 382844 497950 383180 497978
rect 384592 497950 384928 497978
rect 386616 497950 386768 497978
rect 388180 497950 388516 497978
rect 389928 497950 390264 497978
rect 391952 497950 392012 497978
rect 393424 497950 393760 497978
rect 395172 497950 395508 497978
rect 396920 497950 397256 497978
rect 398852 497950 399004 497978
rect 402164 497950 402500 497978
rect 403912 497950 404248 497978
rect 405752 497950 405996 497978
rect 407408 497950 407744 497978
rect 409156 497950 409492 497978
rect 411272 497950 411332 497978
rect 412836 497950 413080 497978
rect 416240 497950 416576 497978
rect 421484 497950 421820 497978
rect 431972 497950 432308 497978
rect 400494 497584 400550 497593
rect 418158 497584 418214 497593
rect 400550 497542 400752 497570
rect 400494 497519 400550 497528
rect 418214 497542 418324 497570
rect 418158 497519 418214 497528
rect 278228 497480 278280 497486
rect 237930 497448 237986 497457
rect 237636 497406 237930 497434
rect 251914 497448 251970 497457
rect 251620 497406 251914 497434
rect 237930 497383 237986 497392
rect 257158 497448 257214 497457
rect 256864 497406 257158 497434
rect 251914 497383 251970 497392
rect 262310 497448 262366 497457
rect 262200 497406 262310 497434
rect 257158 497383 257214 497392
rect 277932 497428 278228 497434
rect 279976 497480 280028 497486
rect 277932 497422 278280 497428
rect 279680 497428 279976 497434
rect 281540 497480 281592 497486
rect 279680 497422 280028 497428
rect 281428 497428 281540 497434
rect 283472 497480 283524 497486
rect 281428 497422 281592 497428
rect 283176 497428 283472 497434
rect 285220 497480 285272 497486
rect 283176 497422 283524 497428
rect 284924 497428 285220 497434
rect 286876 497480 286928 497486
rect 284924 497422 285272 497428
rect 286764 497428 286876 497434
rect 290556 497480 290608 497486
rect 286764 497422 286928 497428
rect 290260 497428 290556 497434
rect 292304 497480 292356 497486
rect 290260 497422 290608 497428
rect 292008 497428 292304 497434
rect 292008 497422 292356 497428
rect 414478 497448 414534 497457
rect 277932 497406 278268 497422
rect 279680 497406 280016 497422
rect 281428 497406 281580 497422
rect 283176 497406 283512 497422
rect 284924 497406 285260 497422
rect 286764 497406 286916 497422
rect 290260 497406 290596 497422
rect 292008 497406 292344 497422
rect 262310 497383 262366 497392
rect 419722 497448 419778 497457
rect 414534 497406 414828 497434
rect 414478 497383 414534 497392
rect 423862 497448 423918 497457
rect 419778 497406 420072 497434
rect 423568 497406 423862 497434
rect 419722 497383 419778 497392
rect 423862 497383 423918 497392
rect 425150 497448 425206 497457
rect 426714 497448 426770 497457
rect 425206 497406 425316 497434
rect 425150 497383 425206 497392
rect 428462 497448 428518 497457
rect 426770 497406 427064 497434
rect 426714 497383 426770 497392
rect 430210 497448 430266 497457
rect 428518 497406 428812 497434
rect 428462 497383 428518 497392
rect 433706 497448 433762 497457
rect 430266 497406 430560 497434
rect 430210 497383 430266 497392
rect 433762 497406 434056 497434
rect 433706 497383 433762 497392
rect 235078 496088 235134 496097
rect 235078 496023 235134 496032
rect 235092 338298 235120 496023
rect 235080 338292 235132 338298
rect 235080 338234 235132 338240
rect 234632 338150 235244 338178
rect 314856 338150 315100 338178
rect 234528 255264 234580 255270
rect 234528 255206 234580 255212
rect 234436 241460 234488 241466
rect 234436 241402 234488 241408
rect 234344 215280 234396 215286
rect 234344 215222 234396 215228
rect 234252 202836 234304 202842
rect 234252 202778 234304 202784
rect 234160 189032 234212 189038
rect 234160 188974 234212 188980
rect 234068 164212 234120 164218
rect 234068 164154 234120 164160
rect 233976 137964 234028 137970
rect 233976 137906 234028 137912
rect 233884 111784 233936 111790
rect 233884 111726 233936 111732
rect 191840 18556 191892 18562
rect 191840 18498 191892 18504
rect 191852 16574 191880 18498
rect 194600 18488 194652 18494
rect 194600 18430 194652 18436
rect 194612 16574 194640 18430
rect 198740 18420 198792 18426
rect 198740 18362 198792 18368
rect 197360 17740 197412 17746
rect 197360 17682 197412 17688
rect 197372 16574 197400 17682
rect 191852 16546 192064 16574
rect 194612 16546 195192 16574
rect 197372 16546 197952 16574
rect 190828 7472 190880 7478
rect 190828 7414 190880 7420
rect 188344 5160 188396 5166
rect 188344 5102 188396 5108
rect 189724 5160 189776 5166
rect 189724 5102 189776 5108
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 189736 480 189764 5102
rect 190840 480 190868 7414
rect 192036 480 192064 16546
rect 194416 7404 194468 7410
rect 194416 7346 194468 7352
rect 193220 5228 193272 5234
rect 193220 5170 193272 5176
rect 193232 480 193260 5170
rect 194428 480 194456 7346
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196808 5296 196860 5302
rect 196808 5238 196860 5244
rect 196820 480 196848 5238
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 18362
rect 208400 17944 208452 17950
rect 208400 17886 208452 17892
rect 204260 17876 204312 17882
rect 204260 17818 204312 17824
rect 201500 17808 201552 17814
rect 201500 17750 201552 17756
rect 200302 4856 200358 4865
rect 200302 4791 200358 4800
rect 200316 480 200344 4791
rect 201512 480 201540 17750
rect 204272 16574 204300 17818
rect 208412 16574 208440 17886
rect 211160 17196 211212 17202
rect 211160 17138 211212 17144
rect 211172 16574 211200 17138
rect 224960 17128 225012 17134
rect 224960 17070 225012 17076
rect 224972 16574 225000 17070
rect 227720 17060 227772 17066
rect 227720 17002 227772 17008
rect 227732 16574 227760 17002
rect 204272 16546 205128 16574
rect 208412 16546 208624 16574
rect 211172 16546 211752 16574
rect 224972 16546 225184 16574
rect 227732 16546 228312 16574
rect 202696 12096 202748 12102
rect 202696 12038 202748 12044
rect 202708 480 202736 12038
rect 203892 5364 203944 5370
rect 203892 5306 203944 5312
rect 203904 480 203932 5306
rect 205100 480 205128 16546
rect 206192 12164 206244 12170
rect 206192 12106 206244 12112
rect 206204 480 206232 12106
rect 207388 5432 207440 5438
rect 207388 5374 207440 5380
rect 207400 480 207428 5374
rect 208596 480 208624 16546
rect 209780 12232 209832 12238
rect 209780 12174 209832 12180
rect 209792 480 209820 12174
rect 210976 5500 211028 5506
rect 210976 5442 211028 5448
rect 210988 480 211016 5442
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 221096 15700 221148 15706
rect 221096 15642 221148 15648
rect 219992 12436 220044 12442
rect 219992 12378 220044 12384
rect 216864 12368 216916 12374
rect 216864 12310 216916 12316
rect 213368 12300 213420 12306
rect 213368 12242 213420 12248
rect 213380 480 213408 12242
rect 215668 9512 215720 9518
rect 215668 9454 215720 9460
rect 214472 4752 214524 4758
rect 214472 4694 214524 4700
rect 214484 480 214512 4694
rect 215680 480 215708 9454
rect 216876 480 216904 12310
rect 219256 9580 219308 9586
rect 219256 9522 219308 9528
rect 218060 4684 218112 4690
rect 218060 4626 218112 4632
rect 218072 480 218100 4626
rect 219268 480 219296 9522
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 12378
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 15642
rect 223580 11688 223632 11694
rect 223580 11630 223632 11636
rect 222752 9648 222804 9654
rect 222752 9590 222804 9596
rect 222764 480 222792 9590
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 11630
rect 225156 480 225184 16546
rect 226340 11620 226392 11626
rect 226340 11562 226392 11568
rect 226352 4214 226380 11562
rect 226432 8900 226484 8906
rect 226432 8842 226484 8848
rect 226340 4208 226392 4214
rect 226340 4150 226392 4156
rect 226444 3482 226472 8842
rect 227536 4208 227588 4214
rect 227536 4150 227588 4156
rect 226352 3454 226472 3482
rect 226352 480 226380 3454
rect 227548 480 227576 4150
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 231032 11552 231084 11558
rect 231032 11494 231084 11500
rect 229836 8832 229888 8838
rect 229836 8774 229888 8780
rect 229848 480 229876 8774
rect 231044 480 231072 11494
rect 233424 8764 233476 8770
rect 233424 8706 233476 8712
rect 232226 6216 232282 6225
rect 232226 6151 232282 6160
rect 232240 480 232268 6151
rect 233436 480 233464 8706
rect 234632 6186 234660 338150
rect 235080 338020 235132 338026
rect 235080 337962 235132 337968
rect 235368 338014 235612 338042
rect 235736 338014 235980 338042
rect 236104 338014 236440 338042
rect 236564 338014 236808 338042
rect 236932 338014 237268 338042
rect 237392 338014 237636 338042
rect 237760 338014 238004 338042
rect 238128 338014 238464 338042
rect 234804 330540 234856 330546
rect 234804 330482 234856 330488
rect 234712 330472 234764 330478
rect 234712 330414 234764 330420
rect 234724 6322 234752 330414
rect 234712 6316 234764 6322
rect 234712 6258 234764 6264
rect 234816 6254 234844 330482
rect 235092 150414 235120 337962
rect 235368 330546 235396 338014
rect 235356 330540 235408 330546
rect 235356 330482 235408 330488
rect 235736 330478 235764 338014
rect 235724 330472 235776 330478
rect 235724 330414 235776 330420
rect 235080 150408 235132 150414
rect 235080 150350 235132 150356
rect 236104 8974 236132 338014
rect 236564 316034 236592 338014
rect 236932 336054 236960 338014
rect 236920 336048 236972 336054
rect 236920 335990 236972 335996
rect 236644 335776 236696 335782
rect 236644 335718 236696 335724
rect 236196 316006 236592 316034
rect 236092 8968 236144 8974
rect 236092 8910 236144 8916
rect 234804 6248 234856 6254
rect 234804 6190 234856 6196
rect 235816 6248 235868 6254
rect 235816 6190 235868 6196
rect 234620 6180 234672 6186
rect 234620 6122 234672 6128
rect 234620 5908 234672 5914
rect 234620 5850 234672 5856
rect 234632 480 234660 5850
rect 235828 480 235856 6190
rect 236196 3369 236224 316006
rect 236182 3360 236238 3369
rect 236182 3295 236238 3304
rect 236656 3262 236684 335718
rect 237392 6390 237420 338014
rect 237760 335354 237788 338014
rect 237484 335326 237788 335354
rect 237484 9042 237512 335326
rect 238128 316034 238156 338014
rect 238818 337770 238846 338028
rect 238956 338014 239292 338042
rect 239416 338014 239660 338042
rect 239784 338014 240028 338042
rect 240152 338014 240488 338042
rect 240612 338014 240856 338042
rect 240980 338014 241316 338042
rect 241532 338014 241684 338042
rect 241808 338014 242052 338042
rect 242176 338014 242512 338042
rect 242636 338014 242880 338042
rect 243096 338014 243340 338042
rect 243464 338014 243708 338042
rect 243832 338014 244168 338042
rect 244476 338014 244536 338042
rect 244660 338014 244904 338042
rect 245028 338014 245364 338042
rect 238818 337742 238892 337770
rect 238760 330540 238812 330546
rect 238760 330482 238812 330488
rect 237576 316006 238156 316034
rect 237576 18601 237604 316006
rect 237562 18592 237618 18601
rect 237562 18527 237618 18536
rect 237472 9036 237524 9042
rect 237472 8978 237524 8984
rect 238116 8968 238168 8974
rect 238116 8910 238168 8916
rect 237380 6384 237432 6390
rect 237380 6326 237432 6332
rect 237012 6180 237064 6186
rect 237012 6122 237064 6128
rect 236644 3256 236696 3262
rect 236644 3198 236696 3204
rect 237024 480 237052 6122
rect 238128 480 238156 8910
rect 238772 3534 238800 330482
rect 238760 3528 238812 3534
rect 238760 3470 238812 3476
rect 238864 3466 238892 337742
rect 238956 6458 238984 338014
rect 239416 316034 239444 338014
rect 239784 330546 239812 338014
rect 240152 336122 240180 338014
rect 240140 336116 240192 336122
rect 240140 336058 240192 336064
rect 239772 330540 239824 330546
rect 239772 330482 239824 330488
rect 240232 330540 240284 330546
rect 240232 330482 240284 330488
rect 239048 316006 239444 316034
rect 239048 11665 239076 316006
rect 240244 13025 240272 330482
rect 240612 316034 240640 338014
rect 240980 330546 241008 338014
rect 240968 330540 241020 330546
rect 240968 330482 241020 330488
rect 240336 316006 240640 316034
rect 240230 13016 240286 13025
rect 240230 12951 240286 12960
rect 239034 11656 239090 11665
rect 239034 11591 239090 11600
rect 240336 6526 240364 316006
rect 240324 6520 240376 6526
rect 240324 6462 240376 6468
rect 238944 6452 238996 6458
rect 238944 6394 238996 6400
rect 239312 6384 239364 6390
rect 239312 6326 239364 6332
rect 238852 3460 238904 3466
rect 238852 3402 238904 3408
rect 239324 480 239352 6326
rect 240508 6316 240560 6322
rect 240508 6258 240560 6264
rect 240520 480 240548 6258
rect 241532 3602 241560 338014
rect 241808 336682 241836 338014
rect 241624 336654 241836 336682
rect 241624 3670 241652 336654
rect 242176 335354 242204 338014
rect 241716 335326 242204 335354
rect 241716 9110 241744 335326
rect 242636 316034 242664 338014
rect 242992 326256 243044 326262
rect 242992 326198 243044 326204
rect 241808 316006 242664 316034
rect 241808 14521 241836 316006
rect 241794 14512 241850 14521
rect 241794 14447 241850 14456
rect 243004 9178 243032 326198
rect 242992 9172 243044 9178
rect 242992 9114 243044 9120
rect 241704 9104 241756 9110
rect 241704 9046 241756 9052
rect 242072 9036 242124 9042
rect 242072 8978 242124 8984
rect 241612 3664 241664 3670
rect 241612 3606 241664 3612
rect 241520 3596 241572 3602
rect 241520 3538 241572 3544
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 228702 -960 228814 326
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 354 241786 480
rect 242084 354 242112 8978
rect 243096 3738 243124 338014
rect 243464 336190 243492 338014
rect 243452 336184 243504 336190
rect 243452 336126 243504 336132
rect 243832 326262 243860 338014
rect 244280 330540 244332 330546
rect 244280 330482 244332 330488
rect 243820 326256 243872 326262
rect 243820 326198 243872 326204
rect 244292 3806 244320 330482
rect 244372 330472 244424 330478
rect 244372 330414 244424 330420
rect 244384 9246 244412 330414
rect 244476 15910 244504 338014
rect 244660 330546 244688 338014
rect 244648 330540 244700 330546
rect 244648 330482 244700 330488
rect 245028 330478 245056 338014
rect 245718 337770 245746 338028
rect 245856 338014 246192 338042
rect 246316 338014 246560 338042
rect 246684 338014 246928 338042
rect 247052 338014 247388 338042
rect 247512 338014 247756 338042
rect 247880 338014 248216 338042
rect 248432 338014 248584 338042
rect 248708 338014 248952 338042
rect 249076 338014 249412 338042
rect 249536 338014 249780 338042
rect 249996 338014 250240 338042
rect 250364 338014 250608 338042
rect 250732 338014 250976 338042
rect 251192 338014 251436 338042
rect 251560 338014 251804 338042
rect 251928 338014 252264 338042
rect 245718 337742 245792 337770
rect 245016 330472 245068 330478
rect 245016 330414 245068 330420
rect 245764 15978 245792 337742
rect 245856 336258 245884 338014
rect 245844 336252 245896 336258
rect 245844 336194 245896 336200
rect 245844 330540 245896 330546
rect 245844 330482 245896 330488
rect 245856 16046 245884 330482
rect 246316 316034 246344 338014
rect 246684 330546 246712 338014
rect 246672 330540 246724 330546
rect 246672 330482 246724 330488
rect 245948 316006 246344 316034
rect 245844 16040 245896 16046
rect 245844 15982 245896 15988
rect 245752 15972 245804 15978
rect 245752 15914 245804 15920
rect 244464 15904 244516 15910
rect 244464 15846 244516 15852
rect 245948 9314 245976 316006
rect 245936 9308 245988 9314
rect 245936 9250 245988 9256
rect 244372 9240 244424 9246
rect 244372 9182 244424 9188
rect 247052 3874 247080 338014
rect 247512 335354 247540 338014
rect 247144 335326 247540 335354
rect 247144 9382 247172 335326
rect 247880 316034 247908 338014
rect 248432 336326 248460 338014
rect 248708 336682 248736 338014
rect 248524 336654 248736 336682
rect 248420 336320 248472 336326
rect 248420 336262 248472 336268
rect 247236 316006 247908 316034
rect 247236 18630 247264 316006
rect 247224 18624 247276 18630
rect 247224 18566 247276 18572
rect 248524 13122 248552 336654
rect 249076 335354 249104 338014
rect 248616 335326 249104 335354
rect 248616 18698 248644 335326
rect 249536 316034 249564 338014
rect 249892 330540 249944 330546
rect 249892 330482 249944 330488
rect 248708 316006 249564 316034
rect 248604 18692 248656 18698
rect 248604 18634 248656 18640
rect 248512 13116 248564 13122
rect 248512 13058 248564 13064
rect 247132 9376 247184 9382
rect 247132 9318 247184 9324
rect 248708 3942 248736 316006
rect 249904 18766 249932 330482
rect 249892 18760 249944 18766
rect 249892 18702 249944 18708
rect 249996 13190 250024 338014
rect 250364 330546 250392 338014
rect 250732 336394 250760 338014
rect 250720 336388 250772 336394
rect 250720 336330 250772 336336
rect 250352 330540 250404 330546
rect 250352 330482 250404 330488
rect 249984 13184 250036 13190
rect 249984 13126 250036 13132
rect 251192 6594 251220 338014
rect 251560 335354 251588 338014
rect 251284 335326 251588 335354
rect 251284 13258 251312 335326
rect 251928 316034 251956 338014
rect 252618 337770 252646 338028
rect 252756 338014 253092 338042
rect 253216 338014 253460 338042
rect 253584 338014 253828 338042
rect 254044 338014 254288 338042
rect 254412 338014 254656 338042
rect 254780 338014 255116 338042
rect 255424 338014 255484 338042
rect 255608 338014 255852 338042
rect 255976 338014 256312 338042
rect 256436 338014 256680 338042
rect 256896 338014 257140 338042
rect 257264 338014 257508 338042
rect 257632 338014 257876 338042
rect 258276 338014 258336 338042
rect 258460 338014 258704 338042
rect 258828 338014 259164 338042
rect 259532 338014 259776 338042
rect 252618 337742 252692 337770
rect 252560 330540 252612 330546
rect 252560 330482 252612 330488
rect 251376 316006 251956 316034
rect 251376 18834 251404 316006
rect 251364 18828 251416 18834
rect 251364 18770 251416 18776
rect 251272 13252 251324 13258
rect 251272 13194 251324 13200
rect 252376 9104 252428 9110
rect 252376 9046 252428 9052
rect 251180 6588 251232 6594
rect 251180 6530 251232 6536
rect 251180 6452 251232 6458
rect 251180 6394 251232 6400
rect 248696 3936 248748 3942
rect 248696 3878 248748 3884
rect 247040 3868 247092 3874
rect 247040 3810 247092 3816
rect 248788 3868 248840 3874
rect 248788 3810 248840 3816
rect 244280 3800 244332 3806
rect 244280 3742 244332 3748
rect 245200 3800 245252 3806
rect 245200 3742 245252 3748
rect 243084 3732 243136 3738
rect 243084 3674 243136 3680
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242912 480 242940 3402
rect 244094 3360 244150 3369
rect 244094 3295 244150 3304
rect 244108 480 244136 3295
rect 245212 480 245240 3742
rect 246396 3528 246448 3534
rect 246396 3470 246448 3476
rect 246408 480 246436 3470
rect 247592 3188 247644 3194
rect 247592 3130 247644 3136
rect 247604 480 247632 3130
rect 248800 480 248828 3810
rect 249984 3596 250036 3602
rect 249984 3538 250036 3544
rect 249996 480 250024 3538
rect 251192 480 251220 6394
rect 252388 480 252416 9046
rect 252572 6730 252600 330482
rect 252560 6724 252612 6730
rect 252560 6666 252612 6672
rect 252664 6662 252692 337742
rect 252756 13326 252784 338014
rect 253216 316034 253244 338014
rect 253584 330546 253612 338014
rect 253572 330540 253624 330546
rect 253572 330482 253624 330488
rect 253940 329996 253992 330002
rect 253940 329938 253992 329944
rect 252848 316006 253244 316034
rect 252848 18902 252876 316006
rect 252836 18896 252888 18902
rect 252836 18838 252888 18844
rect 252744 13320 252796 13326
rect 252744 13262 252796 13268
rect 253952 6798 253980 329938
rect 254044 13394 254072 338014
rect 254412 316034 254440 338014
rect 254780 330002 254808 338014
rect 255320 330472 255372 330478
rect 255320 330414 255372 330420
rect 254768 329996 254820 330002
rect 254768 329938 254820 329944
rect 254136 316006 254440 316034
rect 254136 18970 254164 316006
rect 254124 18964 254176 18970
rect 254124 18906 254176 18912
rect 254032 13388 254084 13394
rect 254032 13330 254084 13336
rect 255332 6866 255360 330414
rect 255424 13462 255452 338014
rect 255504 330540 255556 330546
rect 255504 330482 255556 330488
rect 255516 14482 255544 330482
rect 255608 19990 255636 338014
rect 255976 330478 256004 338014
rect 256436 330546 256464 338014
rect 256424 330540 256476 330546
rect 256424 330482 256476 330488
rect 256792 330540 256844 330546
rect 256792 330482 256844 330488
rect 255964 330472 256016 330478
rect 255964 330414 256016 330420
rect 256700 329180 256752 329186
rect 256700 329122 256752 329128
rect 255596 19984 255648 19990
rect 255596 19926 255648 19932
rect 255504 14476 255556 14482
rect 255504 14418 255556 14424
rect 255412 13456 255464 13462
rect 255412 13398 255464 13404
rect 255872 9172 255924 9178
rect 255872 9114 255924 9120
rect 255320 6860 255372 6866
rect 255320 6802 255372 6808
rect 253940 6792 253992 6798
rect 253940 6734 253992 6740
rect 252652 6656 252704 6662
rect 252652 6598 252704 6604
rect 254676 6520 254728 6526
rect 254676 6462 254728 6468
rect 253480 3664 253532 3670
rect 253480 3606 253532 3612
rect 253492 480 253520 3606
rect 254688 480 254716 6462
rect 255884 480 255912 9114
rect 256712 6118 256740 329122
rect 256804 14550 256832 330482
rect 256896 20058 256924 338014
rect 257264 329186 257292 338014
rect 257632 330546 257660 338014
rect 257620 330540 257672 330546
rect 257620 330482 257672 330488
rect 258172 330540 258224 330546
rect 258172 330482 258224 330488
rect 258080 330132 258132 330138
rect 258080 330074 258132 330080
rect 257252 329180 257304 329186
rect 257252 329122 257304 329128
rect 256884 20052 256936 20058
rect 256884 19994 256936 20000
rect 256792 14544 256844 14550
rect 256792 14486 256844 14492
rect 258092 7614 258120 330074
rect 258184 14618 258212 330482
rect 258276 20126 258304 338014
rect 258460 330138 258488 338014
rect 258828 330546 258856 338014
rect 259460 336796 259512 336802
rect 259460 336738 259512 336744
rect 258816 330540 258868 330546
rect 258816 330482 258868 330488
rect 258448 330132 258500 330138
rect 258448 330074 258500 330080
rect 258264 20120 258316 20126
rect 258264 20062 258316 20068
rect 258172 14612 258224 14618
rect 258172 14554 258224 14560
rect 259472 10305 259500 336738
rect 259552 330540 259604 330546
rect 259552 330482 259604 330488
rect 259564 14686 259592 330482
rect 259644 330472 259696 330478
rect 259644 330414 259696 330420
rect 259656 20262 259684 330414
rect 259644 20256 259696 20262
rect 259644 20198 259696 20204
rect 259748 20194 259776 338014
rect 259840 338014 259900 338042
rect 260024 338014 260360 338042
rect 260484 338014 260728 338042
rect 261036 338014 261188 338042
rect 261312 338014 261556 338042
rect 261680 338014 262016 338042
rect 259840 336802 259868 338014
rect 259828 336796 259880 336802
rect 259828 336738 259880 336744
rect 260024 330546 260052 338014
rect 260104 335708 260156 335714
rect 260104 335650 260156 335656
rect 260012 330540 260064 330546
rect 260012 330482 260064 330488
rect 259736 20188 259788 20194
rect 259736 20130 259788 20136
rect 259552 14680 259604 14686
rect 259552 14622 259604 14628
rect 259458 10296 259514 10305
rect 259458 10231 259514 10240
rect 259460 9240 259512 9246
rect 259460 9182 259512 9188
rect 258080 7608 258132 7614
rect 258080 7550 258132 7556
rect 258264 6588 258316 6594
rect 258264 6530 258316 6536
rect 256700 6112 256752 6118
rect 256700 6054 256752 6060
rect 257068 3732 257120 3738
rect 257068 3674 257120 3680
rect 257080 480 257108 3674
rect 258276 480 258304 6530
rect 259472 480 259500 9182
rect 260116 4622 260144 335650
rect 260484 330478 260512 338014
rect 260472 330472 260524 330478
rect 260472 330414 260524 330420
rect 260932 327548 260984 327554
rect 260932 327490 260984 327496
rect 260944 14754 260972 327490
rect 260932 14748 260984 14754
rect 260932 14690 260984 14696
rect 261036 10334 261064 338014
rect 261312 327554 261340 338014
rect 261680 336462 261708 338014
rect 262370 337770 262398 338028
rect 262508 338014 262752 338042
rect 262876 338014 263212 338042
rect 263336 338014 263580 338042
rect 263704 338014 264040 338042
rect 264164 338014 264408 338042
rect 264532 338014 264776 338042
rect 265084 338014 265236 338042
rect 265360 338014 265604 338042
rect 265728 338014 266064 338042
rect 266432 338014 266676 338042
rect 262370 337742 262444 337770
rect 261668 336456 261720 336462
rect 261668 336398 261720 336404
rect 261484 336184 261536 336190
rect 261484 336126 261536 336132
rect 261300 327548 261352 327554
rect 261300 327490 261352 327496
rect 261024 10328 261076 10334
rect 261024 10270 261076 10276
rect 260104 4616 260156 4622
rect 260104 4558 260156 4564
rect 260656 3256 260708 3262
rect 260656 3198 260708 3204
rect 260668 480 260696 3198
rect 261496 3194 261524 336126
rect 262220 330540 262272 330546
rect 262220 330482 262272 330488
rect 261760 6656 261812 6662
rect 261760 6598 261812 6604
rect 261484 3188 261536 3194
rect 261484 3130 261536 3136
rect 261772 480 261800 6598
rect 262232 4010 262260 330482
rect 262312 330472 262364 330478
rect 262312 330414 262364 330420
rect 262324 10470 262352 330414
rect 262312 10464 262364 10470
rect 262312 10406 262364 10412
rect 262416 10402 262444 337742
rect 262508 14822 262536 338014
rect 262876 330546 262904 338014
rect 262956 336388 263008 336394
rect 262956 336330 263008 336336
rect 262864 330540 262916 330546
rect 262864 330482 262916 330488
rect 262968 316034 262996 336330
rect 263336 330478 263364 338014
rect 263324 330472 263376 330478
rect 263324 330414 263376 330420
rect 262876 316006 262996 316034
rect 262496 14816 262548 14822
rect 262496 14758 262548 14764
rect 262404 10396 262456 10402
rect 262404 10338 262456 10344
rect 262876 5914 262904 316006
rect 263704 14890 263732 338014
rect 264164 336818 264192 338014
rect 264072 336790 264192 336818
rect 264072 336530 264100 336790
rect 264532 336682 264560 338014
rect 264164 336654 264560 336682
rect 264060 336524 264112 336530
rect 264060 336466 264112 336472
rect 264164 316034 264192 336654
rect 264244 336320 264296 336326
rect 264244 336262 264296 336268
rect 263796 316006 264192 316034
rect 263692 14884 263744 14890
rect 263692 14826 263744 14832
rect 263796 10538 263824 316006
rect 263784 10532 263836 10538
rect 263784 10474 263836 10480
rect 262956 9308 263008 9314
rect 262956 9250 263008 9256
rect 262864 5908 262916 5914
rect 262864 5850 262916 5856
rect 262220 4004 262272 4010
rect 262220 3946 262272 3952
rect 262968 480 262996 9250
rect 264152 4004 264204 4010
rect 264152 3946 264204 3952
rect 264164 480 264192 3946
rect 264256 3806 264284 336262
rect 265084 14958 265112 338014
rect 265360 336598 265388 338014
rect 265348 336592 265400 336598
rect 265348 336534 265400 336540
rect 265728 316034 265756 338014
rect 266360 336048 266412 336054
rect 266360 335990 266412 335996
rect 265176 316006 265756 316034
rect 265072 14952 265124 14958
rect 265072 14894 265124 14900
rect 265176 10606 265204 316006
rect 265164 10600 265216 10606
rect 265164 10542 265216 10548
rect 265348 6724 265400 6730
rect 265348 6666 265400 6672
rect 264244 3800 264296 3806
rect 264244 3742 264296 3748
rect 265360 480 265388 6666
rect 266372 3482 266400 335990
rect 266648 330818 266676 338014
rect 266740 338014 266800 338042
rect 266924 338014 267260 338042
rect 267384 338014 267628 338042
rect 267844 338014 268088 338042
rect 268212 338014 268456 338042
rect 268580 338014 268916 338042
rect 269224 338014 269284 338042
rect 269408 338014 269652 338042
rect 269776 338014 270112 338042
rect 270236 338014 270480 338042
rect 270696 338014 270940 338042
rect 271064 338014 271308 338042
rect 271432 338014 271676 338042
rect 271984 338014 272136 338042
rect 272260 338014 272504 338042
rect 272628 338014 272964 338042
rect 266636 330812 266688 330818
rect 266636 330754 266688 330760
rect 266740 330562 266768 338014
rect 266924 335354 266952 338014
rect 266464 330534 266768 330562
rect 266832 335326 266952 335354
rect 266464 4078 266492 330534
rect 266832 330426 266860 335326
rect 266912 330812 266964 330818
rect 266912 330754 266964 330760
rect 266556 330398 266860 330426
rect 266556 13530 266584 330398
rect 266924 330290 266952 330754
rect 266648 330262 266952 330290
rect 266648 15026 266676 330262
rect 267384 316034 267412 338014
rect 267844 336666 267872 338014
rect 267832 336660 267884 336666
rect 267832 336602 267884 336608
rect 267832 330540 267884 330546
rect 267832 330482 267884 330488
rect 266740 316006 267412 316034
rect 266740 15094 266768 316006
rect 267844 15162 267872 330482
rect 268212 316034 268240 338014
rect 268580 330546 268608 338014
rect 269120 336116 269172 336122
rect 269120 336058 269172 336064
rect 268568 330540 268620 330546
rect 268568 330482 268620 330488
rect 267936 316006 268240 316034
rect 267832 15156 267884 15162
rect 267832 15098 267884 15104
rect 266728 15088 266780 15094
rect 266728 15030 266780 15036
rect 266636 15020 266688 15026
rect 266636 14962 266688 14968
rect 267936 13598 267964 316006
rect 267924 13592 267976 13598
rect 267924 13534 267976 13540
rect 266544 13524 266596 13530
rect 266544 13466 266596 13472
rect 268844 6792 268896 6798
rect 268844 6734 268896 6740
rect 266452 4072 266504 4078
rect 266452 4014 266504 4020
rect 267740 4072 267792 4078
rect 267740 4014 267792 4020
rect 266372 3454 266584 3482
rect 266556 480 266584 3454
rect 267752 480 267780 4014
rect 268856 480 268884 6734
rect 269132 3482 269160 336058
rect 269224 4146 269252 338014
rect 269408 335354 269436 338014
rect 269316 335326 269436 335354
rect 269316 13666 269344 335326
rect 269776 316034 269804 338014
rect 270236 336734 270264 338014
rect 270224 336728 270276 336734
rect 270224 336670 270276 336676
rect 270592 330540 270644 330546
rect 270592 330482 270644 330488
rect 269408 316006 269804 316034
rect 269408 14414 269436 316006
rect 269396 14408 269448 14414
rect 269396 14350 269448 14356
rect 270604 14346 270632 330482
rect 270592 14340 270644 14346
rect 270592 14282 270644 14288
rect 270696 13734 270724 338014
rect 271064 330546 271092 338014
rect 271432 335986 271460 338014
rect 271420 335980 271472 335986
rect 271420 335922 271472 335928
rect 271052 330540 271104 330546
rect 271052 330482 271104 330488
rect 271880 330540 271932 330546
rect 271880 330482 271932 330488
rect 270684 13728 270736 13734
rect 270684 13670 270736 13676
rect 269304 13660 269356 13666
rect 269304 13602 269356 13608
rect 271236 6860 271288 6866
rect 271236 6802 271288 6808
rect 269212 4140 269264 4146
rect 269212 4082 269264 4088
rect 269132 3454 270080 3482
rect 270052 480 270080 3454
rect 271248 480 271276 6802
rect 271892 3398 271920 330482
rect 271984 13802 272012 338014
rect 272260 316034 272288 338014
rect 272628 330546 272656 338014
rect 273318 337770 273346 338028
rect 273456 338014 273700 338042
rect 273824 338014 274160 338042
rect 274284 338014 274528 338042
rect 274744 338014 274988 338042
rect 275112 338014 275356 338042
rect 275480 338014 275724 338042
rect 276184 338014 276336 338042
rect 273318 337742 273392 337770
rect 272616 330540 272668 330546
rect 272616 330482 272668 330488
rect 272076 316006 272288 316034
rect 272076 14278 272104 316006
rect 272064 14272 272116 14278
rect 272064 14214 272116 14220
rect 271972 13796 272024 13802
rect 271972 13738 272024 13744
rect 273364 13054 273392 337742
rect 273456 16114 273484 338014
rect 273628 336252 273680 336258
rect 273628 336194 273680 336200
rect 273536 330540 273588 330546
rect 273536 330482 273588 330488
rect 273548 19038 273576 330482
rect 273536 19032 273588 19038
rect 273536 18974 273588 18980
rect 273444 16108 273496 16114
rect 273444 16050 273496 16056
rect 273352 13048 273404 13054
rect 273352 12990 273404 12996
rect 272432 7608 272484 7614
rect 272432 7550 272484 7556
rect 271880 3392 271932 3398
rect 271880 3334 271932 3340
rect 272444 480 272472 7550
rect 273640 480 273668 336194
rect 273824 335918 273852 338014
rect 273812 335912 273864 335918
rect 273812 335854 273864 335860
rect 274284 330546 274312 338014
rect 274640 336728 274692 336734
rect 274640 336670 274692 336676
rect 274272 330540 274324 330546
rect 274272 330482 274324 330488
rect 274652 3330 274680 336670
rect 274744 16182 274772 338014
rect 275112 336734 275140 338014
rect 275100 336728 275152 336734
rect 275100 336670 275152 336676
rect 275480 316034 275508 338014
rect 276204 330540 276256 330546
rect 276204 330482 276256 330488
rect 276112 330472 276164 330478
rect 276112 330414 276164 330420
rect 274836 316006 275508 316034
rect 274836 19106 274864 316006
rect 274824 19100 274876 19106
rect 274824 19042 274876 19048
rect 276124 16318 276152 330414
rect 276216 19174 276244 330482
rect 276204 19168 276256 19174
rect 276204 19110 276256 19116
rect 276112 16312 276164 16318
rect 276112 16254 276164 16260
rect 276308 16250 276336 338014
rect 276400 338014 276552 338042
rect 276676 338014 277012 338042
rect 277136 338014 277380 338042
rect 277596 338014 277840 338042
rect 277964 338014 278208 338042
rect 278332 338014 278576 338042
rect 278884 338014 279036 338042
rect 279160 338014 279404 338042
rect 279528 338014 279864 338042
rect 280232 338014 280384 338042
rect 276400 335850 276428 338014
rect 276388 335844 276440 335850
rect 276388 335786 276440 335792
rect 276676 330546 276704 338014
rect 276664 330540 276716 330546
rect 276664 330482 276716 330488
rect 277136 330478 277164 338014
rect 277596 335782 277624 338014
rect 277584 335776 277636 335782
rect 277584 335718 277636 335724
rect 277964 335354 277992 338014
rect 277504 335326 277992 335354
rect 277124 330472 277176 330478
rect 277124 330414 277176 330420
rect 277504 16386 277532 335326
rect 278332 316034 278360 338014
rect 278780 330540 278832 330546
rect 278780 330482 278832 330488
rect 277596 316006 278360 316034
rect 277492 16380 277544 16386
rect 277492 16322 277544 16328
rect 276296 16244 276348 16250
rect 276296 16186 276348 16192
rect 274732 16176 274784 16182
rect 274732 16118 274784 16124
rect 277124 9376 277176 9382
rect 277124 9318 277176 9324
rect 274824 4140 274876 4146
rect 274824 4082 274876 4088
rect 274640 3324 274692 3330
rect 274640 3266 274692 3272
rect 274836 480 274864 4082
rect 276020 3936 276072 3942
rect 276020 3878 276072 3884
rect 276032 480 276060 3878
rect 277136 480 277164 9318
rect 277596 7750 277624 316006
rect 277584 7744 277636 7750
rect 277584 7686 277636 7692
rect 278792 4826 278820 330482
rect 278884 7682 278912 338014
rect 279160 330546 279188 338014
rect 279148 330540 279200 330546
rect 279148 330482 279200 330488
rect 279528 316034 279556 338014
rect 280356 330562 280384 338014
rect 280540 338014 280600 338042
rect 280724 338014 281060 338042
rect 281184 338014 281428 338042
rect 281552 338014 281888 338042
rect 282012 338014 282256 338042
rect 282380 338014 282624 338042
rect 282932 338014 283084 338042
rect 283208 338014 283452 338042
rect 283576 338014 283912 338042
rect 284036 338014 284280 338042
rect 284588 338014 284648 338042
rect 284772 338014 285108 338042
rect 285232 338014 285476 338042
rect 285876 338014 285936 338042
rect 286060 338014 286304 338042
rect 286428 338014 286764 338042
rect 287132 338014 287376 338042
rect 280252 330540 280304 330546
rect 280356 330534 280476 330562
rect 280252 330482 280304 330488
rect 280160 326732 280212 326738
rect 280160 326674 280212 326680
rect 278976 316006 279556 316034
rect 278976 7818 279004 316006
rect 278964 7812 279016 7818
rect 278964 7754 279016 7760
rect 278872 7676 278924 7682
rect 278872 7618 278924 7624
rect 279516 7676 279568 7682
rect 279516 7618 279568 7624
rect 278780 4820 278832 4826
rect 278780 4762 278832 4768
rect 278320 3392 278372 3398
rect 278320 3334 278372 3340
rect 278332 480 278360 3334
rect 279528 480 279556 7618
rect 280172 4894 280200 326674
rect 280264 8945 280292 330482
rect 280344 330472 280396 330478
rect 280344 330414 280396 330420
rect 280356 11830 280384 330414
rect 280344 11824 280396 11830
rect 280344 11766 280396 11772
rect 280448 11762 280476 330534
rect 280540 326738 280568 338014
rect 280724 330546 280752 338014
rect 280712 330540 280764 330546
rect 280712 330482 280764 330488
rect 281184 330478 281212 338014
rect 281172 330472 281224 330478
rect 281172 330414 281224 330420
rect 280528 326732 280580 326738
rect 280528 326674 280580 326680
rect 280436 11756 280488 11762
rect 280436 11698 280488 11704
rect 280250 8936 280306 8945
rect 280250 8871 280306 8880
rect 281552 6050 281580 338014
rect 282012 335354 282040 338014
rect 281644 335326 282040 335354
rect 281644 9450 281672 335326
rect 282380 316034 282408 338014
rect 281736 316006 282408 316034
rect 281736 11898 281764 316006
rect 281724 11892 281776 11898
rect 281724 11834 281776 11840
rect 281632 9444 281684 9450
rect 281632 9386 281684 9392
rect 281540 6044 281592 6050
rect 281540 5986 281592 5992
rect 282932 5982 282960 338014
rect 283012 330540 283064 330546
rect 283012 330482 283064 330488
rect 283024 11966 283052 330482
rect 283104 328500 283156 328506
rect 283104 328442 283156 328448
rect 283116 16454 283144 328442
rect 283208 17241 283236 338014
rect 283576 330546 283604 338014
rect 283564 330540 283616 330546
rect 283564 330482 283616 330488
rect 284036 328506 284064 338014
rect 284300 336456 284352 336462
rect 284300 336398 284352 336404
rect 284024 328500 284076 328506
rect 284024 328442 284076 328448
rect 283194 17232 283250 17241
rect 283194 17167 283250 17176
rect 283104 16448 283156 16454
rect 283104 16390 283156 16396
rect 283012 11960 283064 11966
rect 283012 11902 283064 11908
rect 283104 7744 283156 7750
rect 283104 7686 283156 7692
rect 282920 5976 282972 5982
rect 282920 5918 282972 5924
rect 280160 4888 280212 4894
rect 280160 4830 280212 4836
rect 281908 4820 281960 4826
rect 281908 4762 281960 4768
rect 280712 3800 280764 3806
rect 280712 3742 280764 3748
rect 280724 480 280752 3742
rect 281920 480 281948 4762
rect 283116 480 283144 7686
rect 284312 480 284340 336398
rect 284392 330540 284444 330546
rect 284392 330482 284444 330488
rect 284404 12034 284432 330482
rect 284484 330472 284536 330478
rect 284484 330414 284536 330420
rect 284496 17406 284524 330414
rect 284484 17400 284536 17406
rect 284484 17342 284536 17348
rect 284588 17270 284616 338014
rect 284772 330546 284800 338014
rect 284760 330540 284812 330546
rect 284760 330482 284812 330488
rect 285232 330478 285260 338014
rect 285772 330540 285824 330546
rect 285772 330482 285824 330488
rect 285220 330472 285272 330478
rect 285220 330414 285272 330420
rect 285680 326868 285732 326874
rect 285680 326810 285732 326816
rect 285692 17610 285720 326810
rect 285680 17604 285732 17610
rect 285680 17546 285732 17552
rect 285784 17474 285812 330482
rect 285772 17468 285824 17474
rect 285772 17410 285824 17416
rect 285876 17338 285904 338014
rect 286060 330546 286088 338014
rect 286048 330540 286100 330546
rect 286048 330482 286100 330488
rect 286428 326874 286456 338014
rect 287060 336524 287112 336530
rect 287060 336466 287112 336472
rect 286416 326868 286468 326874
rect 286416 326810 286468 326816
rect 285864 17332 285916 17338
rect 285864 17274 285916 17280
rect 284576 17264 284628 17270
rect 284576 17206 284628 17212
rect 284392 12028 284444 12034
rect 284392 11970 284444 11976
rect 286600 7812 286652 7818
rect 286600 7754 286652 7760
rect 285404 6112 285456 6118
rect 285404 6054 285456 6060
rect 285416 480 285444 6054
rect 286612 480 286640 7754
rect 287072 6914 287100 336466
rect 287244 330540 287296 330546
rect 287244 330482 287296 330488
rect 287152 330472 287204 330478
rect 287152 330414 287204 330420
rect 287164 10674 287192 330414
rect 287256 17678 287284 330482
rect 287244 17672 287296 17678
rect 287244 17614 287296 17620
rect 287348 17542 287376 338014
rect 287440 338014 287500 338042
rect 287624 338014 287960 338042
rect 288084 338014 288328 338042
rect 288636 338014 288788 338042
rect 288912 338014 289156 338042
rect 289280 338014 289524 338042
rect 287440 19242 287468 338014
rect 287624 330546 287652 338014
rect 287612 330540 287664 330546
rect 287612 330482 287664 330488
rect 288084 330478 288112 338014
rect 288440 330540 288492 330546
rect 288440 330482 288492 330488
rect 288072 330472 288124 330478
rect 288072 330414 288124 330420
rect 287428 19236 287480 19242
rect 287428 19178 287480 19184
rect 287336 17536 287388 17542
rect 287336 17478 287388 17484
rect 287152 10668 287204 10674
rect 287152 10610 287204 10616
rect 288452 7886 288480 330482
rect 288532 330472 288584 330478
rect 288532 330414 288584 330420
rect 288544 10742 288572 330414
rect 288636 12986 288664 338014
rect 288912 330546 288940 338014
rect 288900 330540 288952 330546
rect 288900 330482 288952 330488
rect 289280 330478 289308 338014
rect 289970 337770 289998 338028
rect 290108 338014 290352 338042
rect 290476 338014 290812 338042
rect 290936 338014 291180 338042
rect 291488 338014 291548 338042
rect 291672 338014 292008 338042
rect 292132 338014 292376 338042
rect 292776 338014 292836 338042
rect 292960 338014 293204 338042
rect 293328 338014 293664 338042
rect 294032 338014 294184 338042
rect 289970 337742 290044 337770
rect 289820 330540 289872 330546
rect 289820 330482 289872 330488
rect 289268 330472 289320 330478
rect 289268 330414 289320 330420
rect 288624 12980 288676 12986
rect 288624 12922 288676 12928
rect 288532 10736 288584 10742
rect 288532 10678 288584 10684
rect 289832 7954 289860 330482
rect 289912 327956 289964 327962
rect 289912 327898 289964 327904
rect 289924 10810 289952 327898
rect 290016 12918 290044 337742
rect 290108 16522 290136 338014
rect 290476 330546 290504 338014
rect 290464 330540 290516 330546
rect 290464 330482 290516 330488
rect 290936 327962 290964 338014
rect 291200 336592 291252 336598
rect 291200 336534 291252 336540
rect 290924 327956 290976 327962
rect 290924 327898 290976 327904
rect 290096 16516 290148 16522
rect 290096 16458 290148 16464
rect 290004 12912 290056 12918
rect 290004 12854 290056 12860
rect 289912 10804 289964 10810
rect 289912 10746 289964 10752
rect 289820 7948 289872 7954
rect 289820 7890 289872 7896
rect 290740 7948 290792 7954
rect 290740 7890 290792 7896
rect 288440 7880 288492 7886
rect 288440 7822 288492 7828
rect 288532 7880 288584 7886
rect 288532 7822 288584 7828
rect 287072 6886 287376 6914
rect 241674 326 242112 354
rect 241674 -960 241786 326
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 6886
rect 288544 3942 288572 7822
rect 288992 6044 289044 6050
rect 288992 5986 289044 5992
rect 288532 3936 288584 3942
rect 288532 3878 288584 3884
rect 289004 480 289032 5986
rect 290752 3874 290780 7890
rect 291212 6914 291240 336534
rect 291488 330818 291516 338014
rect 291672 335354 291700 338014
rect 291580 335326 291700 335354
rect 291476 330812 291528 330818
rect 291476 330754 291528 330760
rect 291580 330698 291608 335326
rect 291304 330670 291608 330698
rect 291304 7585 291332 330670
rect 291476 330608 291528 330614
rect 291476 330550 291528 330556
rect 291384 330540 291436 330546
rect 291384 330482 291436 330488
rect 291396 10878 291424 330482
rect 291488 16590 291516 330550
rect 292132 330546 292160 338014
rect 292776 330818 292804 338014
rect 292960 335354 292988 338014
rect 292868 335326 292988 335354
rect 292764 330812 292816 330818
rect 292764 330754 292816 330760
rect 292868 330698 292896 335326
rect 292592 330670 292896 330698
rect 292120 330540 292172 330546
rect 292120 330482 292172 330488
rect 291476 16584 291528 16590
rect 291476 16526 291528 16532
rect 291384 10872 291436 10878
rect 291384 10814 291436 10820
rect 292592 8022 292620 330670
rect 292764 330608 292816 330614
rect 292764 330550 292816 330556
rect 292672 330540 292724 330546
rect 292672 330482 292724 330488
rect 292684 10946 292712 330482
rect 292776 15842 292804 330550
rect 293328 330546 293356 338014
rect 293316 330540 293368 330546
rect 293316 330482 293368 330488
rect 294052 330540 294104 330546
rect 294052 330482 294104 330488
rect 292764 15836 292816 15842
rect 292764 15778 292816 15784
rect 294064 11014 294092 330482
rect 294156 15774 294184 338014
rect 294248 338014 294400 338042
rect 294524 338014 294860 338042
rect 294984 338014 295228 338042
rect 295444 338014 295688 338042
rect 295812 338014 296056 338042
rect 296180 338014 296424 338042
rect 296884 338014 297036 338042
rect 294144 15768 294196 15774
rect 294144 15710 294196 15716
rect 294052 11008 294104 11014
rect 294052 10950 294104 10956
rect 292672 10940 292724 10946
rect 292672 10882 292724 10888
rect 294248 8090 294276 338014
rect 294524 330546 294552 338014
rect 294984 335714 295012 338014
rect 294972 335708 295024 335714
rect 294972 335650 295024 335656
rect 294512 330540 294564 330546
rect 294512 330482 294564 330488
rect 295340 329996 295392 330002
rect 295340 329938 295392 329944
rect 294236 8084 294288 8090
rect 294236 8026 294288 8032
rect 292580 8016 292632 8022
rect 292580 7958 292632 7964
rect 291290 7576 291346 7585
rect 291290 7511 291346 7520
rect 291212 6886 291424 6914
rect 290740 3868 290792 3874
rect 290740 3810 290792 3816
rect 290188 3188 290240 3194
rect 290188 3130 290240 3136
rect 290200 480 290228 3130
rect 291396 480 291424 6886
rect 295352 4962 295380 329938
rect 295444 8158 295472 338014
rect 295812 316034 295840 338014
rect 296180 330002 296208 338014
rect 296718 336016 296774 336025
rect 296718 335951 296774 335960
rect 296168 329996 296220 330002
rect 296168 329938 296220 329944
rect 295536 316006 295840 316034
rect 295536 10266 295564 316006
rect 295524 10260 295576 10266
rect 295524 10202 295576 10208
rect 295432 8152 295484 8158
rect 295432 8094 295484 8100
rect 295340 4956 295392 4962
rect 295340 4898 295392 4904
rect 296076 4956 296128 4962
rect 296076 4898 296128 4904
rect 292580 4888 292632 4894
rect 292580 4830 292632 4836
rect 292592 480 292620 4830
rect 294880 3936 294932 3942
rect 294880 3878 294932 3884
rect 293684 3868 293736 3874
rect 293684 3810 293736 3816
rect 293696 480 293724 3810
rect 294892 480 294920 3878
rect 296088 480 296116 4898
rect 296732 3482 296760 335951
rect 296812 330540 296864 330546
rect 296812 330482 296864 330488
rect 296824 5030 296852 330482
rect 296904 327276 296956 327282
rect 296904 327218 296956 327224
rect 296916 8294 296944 327218
rect 296904 8288 296956 8294
rect 296904 8230 296956 8236
rect 297008 8226 297036 338014
rect 297100 338014 297252 338042
rect 297376 338014 297712 338042
rect 297836 338014 298080 338042
rect 298388 338014 298448 338042
rect 298572 338014 298908 338042
rect 299032 338014 299276 338042
rect 299676 338014 299736 338042
rect 299860 338014 300104 338042
rect 300228 338014 300472 338042
rect 300932 338014 301084 338042
rect 297100 10198 297128 338014
rect 297376 330546 297404 338014
rect 297364 330540 297416 330546
rect 297364 330482 297416 330488
rect 297836 327282 297864 338014
rect 298100 336660 298152 336666
rect 298100 336602 298152 336608
rect 297824 327276 297876 327282
rect 297824 327218 297876 327224
rect 297088 10192 297140 10198
rect 297088 10134 297140 10140
rect 296996 8220 297048 8226
rect 296996 8162 297048 8168
rect 296812 5024 296864 5030
rect 296812 4966 296864 4972
rect 298008 4548 298060 4554
rect 298008 4490 298060 4496
rect 296732 3454 297312 3482
rect 297284 480 297312 3454
rect 298020 3262 298048 4490
rect 298008 3256 298060 3262
rect 298008 3198 298060 3204
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 336602
rect 298192 330540 298244 330546
rect 298192 330482 298244 330488
rect 298204 5098 298232 330482
rect 298284 330472 298336 330478
rect 298284 330414 298336 330420
rect 298296 7546 298324 330414
rect 298388 10130 298416 338014
rect 298572 330546 298600 338014
rect 298560 330540 298612 330546
rect 298560 330482 298612 330488
rect 299032 330478 299060 338014
rect 299572 330540 299624 330546
rect 299572 330482 299624 330488
rect 299020 330472 299072 330478
rect 299020 330414 299072 330420
rect 299480 330132 299532 330138
rect 299480 330074 299532 330080
rect 298376 10124 298428 10130
rect 298376 10066 298428 10072
rect 298284 7540 298336 7546
rect 298284 7482 298336 7488
rect 299492 5166 299520 330074
rect 299584 7478 299612 330482
rect 299676 19310 299704 338014
rect 299860 330138 299888 338014
rect 300228 330546 300256 338014
rect 301056 330818 301084 338014
rect 301148 338014 301300 338042
rect 301424 338014 301760 338042
rect 301884 338014 302128 338042
rect 302252 338014 302588 338042
rect 302712 338014 302956 338042
rect 303080 338014 303324 338042
rect 303724 338014 303784 338042
rect 303908 338014 304152 338042
rect 304276 338014 304612 338042
rect 304736 338014 304980 338042
rect 305288 338014 305348 338042
rect 305472 338014 305808 338042
rect 305932 338014 306176 338042
rect 306576 338014 306636 338042
rect 306760 338014 307004 338042
rect 307128 338014 307372 338042
rect 307832 338014 307984 338042
rect 301044 330812 301096 330818
rect 301044 330754 301096 330760
rect 301148 330698 301176 338014
rect 300872 330670 301176 330698
rect 300216 330540 300268 330546
rect 300216 330482 300268 330488
rect 299848 330132 299900 330138
rect 299848 330074 299900 330080
rect 299664 19304 299716 19310
rect 299664 19246 299716 19252
rect 299572 7472 299624 7478
rect 299572 7414 299624 7420
rect 300872 5234 300900 330670
rect 301044 330608 301096 330614
rect 301044 330550 301096 330556
rect 300952 330540 301004 330546
rect 300952 330482 301004 330488
rect 300964 7410 300992 330482
rect 301056 18562 301084 330550
rect 301424 330546 301452 338014
rect 301412 330540 301464 330546
rect 301412 330482 301464 330488
rect 301884 316034 301912 338014
rect 301148 316006 301912 316034
rect 301044 18556 301096 18562
rect 301044 18498 301096 18504
rect 301148 18494 301176 316006
rect 301136 18488 301188 18494
rect 301136 18430 301188 18436
rect 300952 7404 301004 7410
rect 300952 7346 301004 7352
rect 302252 5302 302280 338014
rect 302712 335354 302740 338014
rect 302344 335326 302740 335354
rect 302344 17746 302372 335326
rect 303080 316034 303108 338014
rect 303620 326460 303672 326466
rect 303620 326402 303672 326408
rect 302436 316006 303108 316034
rect 302436 18426 302464 316006
rect 302424 18420 302476 18426
rect 302424 18362 302476 18368
rect 302332 17740 302384 17746
rect 302332 17682 302384 17688
rect 303632 5370 303660 326402
rect 303620 5364 303672 5370
rect 303620 5306 303672 5312
rect 302240 5296 302292 5302
rect 302240 5238 302292 5244
rect 300860 5228 300912 5234
rect 300860 5170 300912 5176
rect 299480 5160 299532 5166
rect 299480 5102 299532 5108
rect 298192 5092 298244 5098
rect 298192 5034 298244 5040
rect 303160 5092 303212 5098
rect 303160 5034 303212 5040
rect 299664 5024 299716 5030
rect 299664 4966 299716 4972
rect 299296 4616 299348 4622
rect 299296 4558 299348 4564
rect 299308 3398 299336 4558
rect 299388 4480 299440 4486
rect 299388 4422 299440 4428
rect 299400 4010 299428 4422
rect 299388 4004 299440 4010
rect 299388 3946 299440 3952
rect 299296 3392 299348 3398
rect 299296 3334 299348 3340
rect 299676 480 299704 4966
rect 301504 4412 301556 4418
rect 301504 4354 301556 4360
rect 301516 4078 301544 4354
rect 301504 4072 301556 4078
rect 301504 4014 301556 4020
rect 300768 3324 300820 3330
rect 300768 3266 300820 3272
rect 300780 480 300808 3266
rect 301964 3120 302016 3126
rect 301964 3062 302016 3068
rect 301976 480 302004 3062
rect 303172 480 303200 5034
rect 303724 4865 303752 338014
rect 303804 326392 303856 326398
rect 303804 326334 303856 326340
rect 303816 12102 303844 326334
rect 303908 17814 303936 338014
rect 304276 326398 304304 338014
rect 304736 326466 304764 338014
rect 305000 336728 305052 336734
rect 305000 336670 305052 336676
rect 304724 326460 304776 326466
rect 304724 326402 304776 326408
rect 304264 326392 304316 326398
rect 304264 326334 304316 326340
rect 303896 17808 303948 17814
rect 303896 17750 303948 17756
rect 303804 12096 303856 12102
rect 303804 12038 303856 12044
rect 303710 4856 303766 4865
rect 303710 4791 303766 4800
rect 305012 3482 305040 336670
rect 305288 326466 305316 338014
rect 305472 335354 305500 338014
rect 305380 335326 305500 335354
rect 305276 326460 305328 326466
rect 305276 326402 305328 326408
rect 305092 326392 305144 326398
rect 305092 326334 305144 326340
rect 305104 5438 305132 326334
rect 305380 323626 305408 335326
rect 305460 326460 305512 326466
rect 305460 326402 305512 326408
rect 305196 323598 305408 323626
rect 305196 12170 305224 323598
rect 305472 318794 305500 326402
rect 305932 326398 305960 338014
rect 306576 326466 306604 338014
rect 306760 335354 306788 338014
rect 306668 335326 306788 335354
rect 306564 326460 306616 326466
rect 306564 326402 306616 326408
rect 305920 326392 305972 326398
rect 305920 326334 305972 326340
rect 306564 326256 306616 326262
rect 306564 326198 306616 326204
rect 306472 323604 306524 323610
rect 306472 323546 306524 323552
rect 306380 322788 306432 322794
rect 306380 322730 306432 322736
rect 305288 318766 305500 318794
rect 305288 17882 305316 318766
rect 305276 17876 305328 17882
rect 305276 17818 305328 17824
rect 305184 12164 305236 12170
rect 305184 12106 305236 12112
rect 306392 5506 306420 322730
rect 306484 12238 306512 323546
rect 306576 17950 306604 326198
rect 306668 323610 306696 335326
rect 306656 323604 306708 323610
rect 306656 323546 306708 323552
rect 307128 322794 307156 338014
rect 307956 336802 307984 338014
rect 308048 338014 308200 338042
rect 308324 338014 308660 338042
rect 308784 338014 309028 338042
rect 309336 338014 309396 338042
rect 309520 338014 309856 338042
rect 309980 338014 310224 338042
rect 307944 336796 307996 336802
rect 307944 336738 307996 336744
rect 307760 335980 307812 335986
rect 307760 335922 307812 335928
rect 307116 322788 307168 322794
rect 307116 322730 307168 322736
rect 306564 17944 306616 17950
rect 306564 17886 306616 17892
rect 306472 12232 306524 12238
rect 306472 12174 306524 12180
rect 306380 5500 306432 5506
rect 306380 5442 306432 5448
rect 305092 5432 305144 5438
rect 305092 5374 305144 5380
rect 306748 5160 306800 5166
rect 306748 5102 306800 5108
rect 305012 3454 305592 3482
rect 304356 3256 304408 3262
rect 304356 3198 304408 3204
rect 304368 480 304396 3198
rect 305564 480 305592 3454
rect 306760 480 306788 5102
rect 307772 3482 307800 335922
rect 307944 326460 307996 326466
rect 307944 326402 307996 326408
rect 307852 326392 307904 326398
rect 307852 326334 307904 326340
rect 307864 4758 307892 326334
rect 307956 9518 307984 326402
rect 308048 12306 308076 338014
rect 308128 336796 308180 336802
rect 308128 336738 308180 336744
rect 308140 17202 308168 336738
rect 308324 326398 308352 338014
rect 308784 326466 308812 338014
rect 309336 328454 309364 338014
rect 309520 335354 309548 338014
rect 309244 328426 309364 328454
rect 309428 335326 309548 335354
rect 309140 326732 309192 326738
rect 309140 326674 309192 326680
rect 308772 326460 308824 326466
rect 308772 326402 308824 326408
rect 308312 326392 308364 326398
rect 308312 326334 308364 326340
rect 308128 17196 308180 17202
rect 308128 17138 308180 17144
rect 308036 12300 308088 12306
rect 308036 12242 308088 12248
rect 307944 9512 307996 9518
rect 307944 9454 307996 9460
rect 307852 4752 307904 4758
rect 307852 4694 307904 4700
rect 309152 4690 309180 326674
rect 309244 326482 309272 328426
rect 309428 326738 309456 335326
rect 309416 326732 309468 326738
rect 309416 326674 309468 326680
rect 309244 326454 309364 326482
rect 309232 326392 309284 326398
rect 309232 326334 309284 326340
rect 309244 9586 309272 326334
rect 309336 12374 309364 326454
rect 309980 326398 310008 338014
rect 310670 337770 310698 338028
rect 310808 338014 311052 338042
rect 311176 338014 311512 338042
rect 311636 338014 311880 338042
rect 312188 338014 312248 338042
rect 312372 338014 312708 338042
rect 312832 338014 313076 338042
rect 313476 338014 313536 338042
rect 313660 338014 313904 338042
rect 314028 338014 314272 338042
rect 310670 337742 310744 337770
rect 310612 326460 310664 326466
rect 310612 326402 310664 326408
rect 309968 326392 310020 326398
rect 309968 326334 310020 326340
rect 310520 326392 310572 326398
rect 310520 326334 310572 326340
rect 309324 12368 309376 12374
rect 309324 12310 309376 12316
rect 310532 9654 310560 326334
rect 310624 11694 310652 326402
rect 310716 12442 310744 337742
rect 310808 15706 310836 338014
rect 311176 326398 311204 338014
rect 311636 326466 311664 338014
rect 311900 335912 311952 335918
rect 311900 335854 311952 335860
rect 311624 326460 311676 326466
rect 311624 326402 311676 326408
rect 311164 326392 311216 326398
rect 311164 326334 311216 326340
rect 310796 15700 310848 15706
rect 310796 15642 310848 15648
rect 310704 12436 310756 12442
rect 310704 12378 310756 12384
rect 310612 11688 310664 11694
rect 310612 11630 310664 11636
rect 310520 9648 310572 9654
rect 310520 9590 310572 9596
rect 309232 9580 309284 9586
rect 309232 9522 309284 9528
rect 311912 6914 311940 335854
rect 311992 330540 312044 330546
rect 311992 330482 312044 330488
rect 312004 8906 312032 330482
rect 312084 330472 312136 330478
rect 312084 330414 312136 330420
rect 312096 11626 312124 330414
rect 312188 17134 312216 338014
rect 312372 330546 312400 338014
rect 312360 330540 312412 330546
rect 312360 330482 312412 330488
rect 312832 330478 312860 338014
rect 313372 330540 313424 330546
rect 313372 330482 313424 330488
rect 312820 330472 312872 330478
rect 312820 330414 312872 330420
rect 313280 328772 313332 328778
rect 313280 328714 313332 328720
rect 312176 17128 312228 17134
rect 312176 17070 312228 17076
rect 312084 11620 312136 11626
rect 312084 11562 312136 11568
rect 311992 8900 312044 8906
rect 311992 8842 312044 8848
rect 313292 8838 313320 328714
rect 313384 11558 313412 330482
rect 313476 17066 313504 338014
rect 313660 328778 313688 338014
rect 314028 330546 314056 338014
rect 314718 337822 314746 338028
rect 314706 337816 314758 337822
rect 314706 337758 314758 337764
rect 314016 330540 314068 330546
rect 314016 330482 314068 330488
rect 314752 330540 314804 330546
rect 314752 330482 314804 330488
rect 313648 328772 313700 328778
rect 313648 328714 313700 328720
rect 313464 17060 313516 17066
rect 313464 17002 313516 17008
rect 313372 11552 313424 11558
rect 313372 11494 313424 11500
rect 313280 8832 313332 8838
rect 313280 8774 313332 8780
rect 311912 6886 312216 6914
rect 309876 5976 309928 5982
rect 309876 5918 309928 5924
rect 309140 4684 309192 4690
rect 309140 4626 309192 4632
rect 309048 4072 309100 4078
rect 309048 4014 309100 4020
rect 307772 3454 307984 3482
rect 307956 480 307984 3454
rect 309060 480 309088 4014
rect 309888 3194 309916 5918
rect 310244 5228 310296 5234
rect 310244 5170 310296 5176
rect 309876 3188 309928 3194
rect 309876 3130 309928 3136
rect 310256 480 310284 5170
rect 311440 4140 311492 4146
rect 311440 4082 311492 4088
rect 311452 480 311480 4082
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 6886
rect 314764 6254 314792 330482
rect 314856 8770 314884 338150
rect 315224 338014 315560 338042
rect 315684 338014 315928 338042
rect 316144 338014 316296 338042
rect 316420 338014 316756 338042
rect 316880 338014 317124 338042
rect 314936 337816 314988 337822
rect 314936 337758 314988 337764
rect 314844 8764 314896 8770
rect 314844 8706 314896 8712
rect 314752 6248 314804 6254
rect 314948 6225 314976 337758
rect 315224 336394 315252 338014
rect 315212 336388 315264 336394
rect 315212 336330 315264 336336
rect 315684 330546 315712 338014
rect 316040 336388 316092 336394
rect 316040 336330 316092 336336
rect 315672 330540 315724 330546
rect 315672 330482 315724 330488
rect 316052 9674 316080 336330
rect 316144 12050 316172 338014
rect 316224 330540 316276 330546
rect 316224 330482 316276 330488
rect 316236 12170 316264 330482
rect 316420 316034 316448 338014
rect 316880 330546 316908 338014
rect 317570 337770 317598 338028
rect 317708 338014 317952 338042
rect 318076 338014 318320 338042
rect 318444 338014 318780 338042
rect 318904 338014 319148 338042
rect 319272 338014 319608 338042
rect 319732 338014 319976 338042
rect 320376 338014 320436 338042
rect 320560 338014 320804 338042
rect 320928 338014 321172 338042
rect 321632 338014 321784 338042
rect 317570 337742 317644 337770
rect 316868 330540 316920 330546
rect 316868 330482 316920 330488
rect 317420 330540 317472 330546
rect 317420 330482 317472 330488
rect 316328 316006 316448 316034
rect 316328 16574 316356 316006
rect 316328 16546 316448 16574
rect 316224 12164 316276 12170
rect 316224 12106 316276 12112
rect 316144 12022 316356 12050
rect 316132 11960 316184 11966
rect 316132 11902 316184 11908
rect 315960 9646 316080 9674
rect 315960 9518 315988 9646
rect 316040 9580 316092 9586
rect 316040 9522 316092 9528
rect 315948 9512 316000 9518
rect 315948 9454 316000 9460
rect 314752 6190 314804 6196
rect 314934 6216 314990 6225
rect 316052 6186 316080 9522
rect 316144 6390 316172 11902
rect 316328 9586 316356 12022
rect 316316 9580 316368 9586
rect 316316 9522 316368 9528
rect 316224 9512 316276 9518
rect 316224 9454 316276 9460
rect 316132 6384 316184 6390
rect 316132 6326 316184 6332
rect 314934 6151 314990 6160
rect 316040 6180 316092 6186
rect 316040 6122 316092 6128
rect 313832 5296 313884 5302
rect 313832 5238 313884 5244
rect 313844 480 313872 5238
rect 315028 3392 315080 3398
rect 315028 3334 315080 3340
rect 315040 480 315068 3334
rect 316236 480 316264 9454
rect 316420 8974 316448 16546
rect 316408 8968 316460 8974
rect 316408 8910 316460 8916
rect 317328 5364 317380 5370
rect 317328 5306 317380 5312
rect 317340 480 317368 5306
rect 317432 3466 317460 330482
rect 317512 330472 317564 330478
rect 317512 330414 317564 330420
rect 317420 3460 317472 3466
rect 317420 3402 317472 3408
rect 317524 3369 317552 330414
rect 317616 6322 317644 337742
rect 317708 9042 317736 338014
rect 318076 330546 318104 338014
rect 318064 330540 318116 330546
rect 318064 330482 318116 330488
rect 318444 330478 318472 338014
rect 318904 336326 318932 338014
rect 318892 336320 318944 336326
rect 318892 336262 318944 336268
rect 318800 335844 318852 335850
rect 318800 335786 318852 335792
rect 318432 330472 318484 330478
rect 318432 330414 318484 330420
rect 317696 9036 317748 9042
rect 317696 8978 317748 8984
rect 317604 6316 317656 6322
rect 317604 6258 317656 6264
rect 317880 4004 317932 4010
rect 317880 3946 317932 3952
rect 317892 3738 317920 3946
rect 317880 3732 317932 3738
rect 317880 3674 317932 3680
rect 318812 3482 318840 335786
rect 319272 316034 319300 338014
rect 319732 336190 319760 338014
rect 319720 336184 319772 336190
rect 319720 336126 319772 336132
rect 320376 330818 320404 338014
rect 320560 335354 320588 338014
rect 320468 335326 320588 335354
rect 320364 330812 320416 330818
rect 320364 330754 320416 330760
rect 320468 330698 320496 335326
rect 318904 316006 319300 316034
rect 320192 330670 320496 330698
rect 318904 3602 318932 316006
rect 320192 3670 320220 330670
rect 320364 330608 320416 330614
rect 320364 330550 320416 330556
rect 320272 330540 320324 330546
rect 320272 330482 320324 330488
rect 320284 6458 320312 330482
rect 320376 7954 320404 330550
rect 320928 330546 320956 338014
rect 321560 336796 321612 336802
rect 321560 336738 321612 336744
rect 320916 330540 320968 330546
rect 320916 330482 320968 330488
rect 320364 7948 320416 7954
rect 320364 7890 320416 7896
rect 320272 6452 320324 6458
rect 320272 6394 320324 6400
rect 321572 3738 321600 336738
rect 321652 330540 321704 330546
rect 321652 330482 321704 330488
rect 321664 6526 321692 330482
rect 321756 9110 321784 338014
rect 321848 338014 322000 338042
rect 322124 338014 322460 338042
rect 322584 338014 322828 338042
rect 322952 338014 323196 338042
rect 323320 338014 323656 338042
rect 323780 338014 324024 338042
rect 324424 338014 324484 338042
rect 324608 338014 324852 338042
rect 324976 338014 325220 338042
rect 325344 338014 325680 338042
rect 325896 338014 326048 338042
rect 326172 338014 326508 338042
rect 326632 338014 326876 338042
rect 327276 338014 327336 338042
rect 327460 338014 327704 338042
rect 327828 338014 328072 338042
rect 328532 338014 328684 338042
rect 321848 336802 321876 338014
rect 321836 336796 321888 336802
rect 321836 336738 321888 336744
rect 322124 330546 322152 338014
rect 322112 330540 322164 330546
rect 322112 330482 322164 330488
rect 322584 316034 322612 338014
rect 321848 316006 322612 316034
rect 321848 9178 321876 316006
rect 321836 9172 321888 9178
rect 321836 9114 321888 9120
rect 321744 9104 321796 9110
rect 321744 9046 321796 9052
rect 321652 6520 321704 6526
rect 321652 6462 321704 6468
rect 322952 4010 322980 338014
rect 323320 335354 323348 338014
rect 323044 335326 323348 335354
rect 323044 6594 323072 335326
rect 323780 316034 323808 338014
rect 324320 330540 324372 330546
rect 324320 330482 324372 330488
rect 323136 316006 323808 316034
rect 323136 9246 323164 316006
rect 323124 9240 323176 9246
rect 323124 9182 323176 9188
rect 323032 6588 323084 6594
rect 323032 6530 323084 6536
rect 324332 5658 324360 330482
rect 324240 5630 324360 5658
rect 324240 4486 324268 5630
rect 324424 5522 324452 338014
rect 324608 335354 324636 338014
rect 324516 335326 324636 335354
rect 324516 6662 324544 335326
rect 324976 316034 325004 338014
rect 325344 330546 325372 338014
rect 325332 330540 325384 330546
rect 325332 330482 325384 330488
rect 325792 326936 325844 326942
rect 325792 326878 325844 326884
rect 324608 316006 325004 316034
rect 324608 9314 324636 316006
rect 324596 9308 324648 9314
rect 324596 9250 324648 9256
rect 324504 6656 324556 6662
rect 324504 6598 324556 6604
rect 324332 5494 324452 5522
rect 324332 4554 324360 5494
rect 324412 5432 324464 5438
rect 324412 5374 324464 5380
rect 324320 4548 324372 4554
rect 324320 4490 324372 4496
rect 324228 4480 324280 4486
rect 324228 4422 324280 4428
rect 322940 4004 322992 4010
rect 322940 3946 322992 3952
rect 321560 3732 321612 3738
rect 321560 3674 321612 3680
rect 320180 3664 320232 3670
rect 320180 3606 320232 3612
rect 318892 3596 318944 3602
rect 318892 3538 318944 3544
rect 323308 3596 323360 3602
rect 323308 3538 323360 3544
rect 322112 3528 322164 3534
rect 318812 3454 319760 3482
rect 322112 3470 322164 3476
rect 317510 3360 317566 3369
rect 317510 3295 317566 3304
rect 318524 3052 318576 3058
rect 318524 2994 318576 3000
rect 318536 480 318564 2994
rect 319732 480 319760 3454
rect 320916 3188 320968 3194
rect 320916 3130 320968 3136
rect 320928 480 320956 3130
rect 322124 480 322152 3470
rect 323320 480 323348 3538
rect 324424 480 324452 5374
rect 325804 4418 325832 326878
rect 325896 6730 325924 338014
rect 326172 336054 326200 338014
rect 326160 336048 326212 336054
rect 326160 335990 326212 335996
rect 326344 335776 326396 335782
rect 326344 335718 326396 335724
rect 325976 335708 326028 335714
rect 325976 335650 326028 335656
rect 325988 6914 326016 335650
rect 326356 16574 326384 335718
rect 326632 326942 326660 338014
rect 327172 330540 327224 330546
rect 327172 330482 327224 330488
rect 326620 326936 326672 326942
rect 326620 326878 326672 326884
rect 326356 16546 326476 16574
rect 325988 6886 326384 6914
rect 325884 6724 325936 6730
rect 325884 6666 325936 6672
rect 325792 4412 325844 4418
rect 325792 4354 325844 4360
rect 325608 3664 325660 3670
rect 325608 3606 325660 3612
rect 325620 480 325648 3606
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 6886
rect 326448 3330 326476 16546
rect 327184 6866 327212 330482
rect 327172 6860 327224 6866
rect 327172 6802 327224 6808
rect 327276 6798 327304 338014
rect 327356 336184 327408 336190
rect 327356 336126 327408 336132
rect 327368 16574 327396 336126
rect 327460 336122 327488 338014
rect 327448 336116 327500 336122
rect 327448 336058 327500 336064
rect 327828 330546 327856 338014
rect 327816 330540 327868 330546
rect 327816 330482 327868 330488
rect 328552 330540 328604 330546
rect 328552 330482 328604 330488
rect 327368 16546 328040 16574
rect 327264 6792 327316 6798
rect 327264 6734 327316 6740
rect 326436 3324 326488 3330
rect 326436 3266 326488 3272
rect 328012 480 328040 16546
rect 328564 7886 328592 330482
rect 328552 7880 328604 7886
rect 328552 7822 328604 7828
rect 328656 7614 328684 338014
rect 328748 338014 328900 338042
rect 329024 338014 329360 338042
rect 329484 338014 329728 338042
rect 330036 338014 330096 338042
rect 330220 338014 330556 338042
rect 330680 338014 330924 338042
rect 331324 338014 331384 338042
rect 331508 338014 331752 338042
rect 331876 338014 332120 338042
rect 332244 338014 332580 338042
rect 332796 338014 332948 338042
rect 333072 338014 333408 338042
rect 333532 338014 333776 338042
rect 334084 338014 334144 338042
rect 334268 338014 334604 338042
rect 334728 338014 334972 338042
rect 335432 338014 335584 338042
rect 328748 336258 328776 338014
rect 328920 336592 328972 336598
rect 328920 336534 328972 336540
rect 328932 336326 328960 336534
rect 328920 336320 328972 336326
rect 328920 336262 328972 336268
rect 328736 336252 328788 336258
rect 328736 336194 328788 336200
rect 329024 316034 329052 338014
rect 329104 335640 329156 335646
rect 329104 335582 329156 335588
rect 328748 316006 329052 316034
rect 328644 7608 328696 7614
rect 328644 7550 328696 7556
rect 328748 4350 328776 316006
rect 328736 4344 328788 4350
rect 328736 4286 328788 4292
rect 329116 3262 329144 335582
rect 329484 330546 329512 338014
rect 329472 330540 329524 330546
rect 329472 330482 329524 330488
rect 329840 327820 329892 327826
rect 329840 327762 329892 327768
rect 329852 4622 329880 327762
rect 329932 326868 329984 326874
rect 329932 326810 329984 326816
rect 329944 7682 329972 326810
rect 330036 9382 330064 338014
rect 330220 327826 330248 338014
rect 330208 327820 330260 327826
rect 330208 327762 330260 327768
rect 330680 326874 330708 338014
rect 331220 336048 331272 336054
rect 331220 335990 331272 335996
rect 330668 326868 330720 326874
rect 330668 326810 330720 326816
rect 330024 9376 330076 9382
rect 330024 9318 330076 9324
rect 329932 7676 329984 7682
rect 329932 7618 329984 7624
rect 329840 4616 329892 4622
rect 329840 4558 329892 4564
rect 330392 3732 330444 3738
rect 330392 3674 330444 3680
rect 329196 3460 329248 3466
rect 329196 3402 329248 3408
rect 329104 3256 329156 3262
rect 329104 3198 329156 3204
rect 329208 480 329236 3402
rect 330404 480 330432 3674
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 335990
rect 331324 3806 331352 338014
rect 331508 335354 331536 338014
rect 331876 336682 331904 338014
rect 331416 335326 331536 335354
rect 331784 336654 331904 336682
rect 331416 4826 331444 335326
rect 331784 316034 331812 336654
rect 332244 336530 332272 338014
rect 332232 336524 332284 336530
rect 332232 336466 332284 336472
rect 331864 336456 331916 336462
rect 331864 336398 331916 336404
rect 331508 316006 331812 316034
rect 331508 7750 331536 316006
rect 331496 7744 331548 7750
rect 331496 7686 331548 7692
rect 331404 4820 331456 4826
rect 331404 4762 331456 4768
rect 331312 3800 331364 3806
rect 331312 3742 331364 3748
rect 331876 3194 331904 336398
rect 332692 326392 332744 326398
rect 332692 326334 332744 326340
rect 332704 7818 332732 326334
rect 332692 7812 332744 7818
rect 332692 7754 332744 7760
rect 332796 6118 332824 338014
rect 333072 326398 333100 338014
rect 333532 336598 333560 338014
rect 333520 336592 333572 336598
rect 333520 336534 333572 336540
rect 333244 335572 333296 335578
rect 333244 335514 333296 335520
rect 333060 326392 333112 326398
rect 333060 326334 333112 326340
rect 332784 6112 332836 6118
rect 332784 6054 332836 6060
rect 332692 3800 332744 3806
rect 332692 3742 332744 3748
rect 331864 3188 331916 3194
rect 331864 3130 331916 3136
rect 332704 480 332732 3742
rect 333256 3466 333284 335514
rect 334084 6050 334112 338014
rect 334268 316034 334296 338014
rect 334728 336326 334756 338014
rect 334716 336320 334768 336326
rect 334716 336262 334768 336268
rect 334992 336252 335044 336258
rect 334992 336194 335044 336200
rect 334900 336184 334952 336190
rect 334900 336126 334952 336132
rect 334624 336116 334676 336122
rect 334624 336058 334676 336064
rect 334176 316006 334296 316034
rect 334072 6044 334124 6050
rect 334072 5986 334124 5992
rect 334176 5982 334204 316006
rect 334164 5976 334216 5982
rect 334164 5918 334216 5924
rect 334636 3466 334664 336058
rect 334912 335714 334940 336126
rect 334900 335708 334952 335714
rect 334900 335650 334952 335656
rect 335004 335578 335032 336194
rect 334992 335572 335044 335578
rect 334992 335514 335044 335520
rect 335556 326466 335584 338014
rect 335740 338014 335800 338042
rect 335924 338014 336260 338042
rect 336384 338014 336628 338042
rect 336752 338014 336996 338042
rect 337120 338014 337456 338042
rect 337580 338014 337824 338042
rect 338132 338014 338284 338042
rect 338408 338014 338652 338042
rect 338776 338014 339020 338042
rect 339144 338014 339480 338042
rect 339604 338014 339848 338042
rect 339972 338014 340308 338042
rect 340432 338014 340676 338042
rect 340892 338014 341044 338042
rect 341168 338014 341504 338042
rect 341628 338014 341872 338042
rect 342272 338014 342332 338042
rect 342456 338014 342700 338042
rect 342824 338014 343068 338042
rect 343192 338014 343528 338042
rect 343744 338014 343896 338042
rect 344020 338014 344356 338042
rect 344480 338014 344724 338042
rect 345032 338014 345184 338042
rect 345308 338014 345552 338042
rect 345676 338014 345920 338042
rect 346044 338014 346380 338042
rect 346504 338014 346748 338042
rect 346872 338014 347208 338042
rect 347332 338014 347576 338042
rect 347792 338014 347944 338042
rect 348068 338014 348404 338042
rect 348528 338014 348772 338042
rect 349232 338014 349476 338042
rect 335544 326460 335596 326466
rect 335544 326402 335596 326408
rect 335360 326392 335412 326398
rect 335740 326346 335768 338014
rect 335820 326460 335872 326466
rect 335820 326402 335872 326408
rect 335360 326334 335412 326340
rect 335372 3942 335400 326334
rect 335464 326318 335768 326346
rect 335360 3936 335412 3942
rect 335360 3878 335412 3884
rect 335464 3874 335492 326318
rect 335544 326256 335596 326262
rect 335544 326198 335596 326204
rect 335556 4962 335584 326198
rect 335832 321554 335860 326402
rect 335924 326398 335952 338014
rect 335912 326392 335964 326398
rect 335912 326334 335964 326340
rect 336384 326262 336412 338014
rect 336752 336025 336780 338014
rect 337120 336666 337148 338014
rect 337108 336660 337160 336666
rect 337108 336602 337160 336608
rect 336738 336016 336794 336025
rect 336738 335951 336794 335960
rect 336372 326256 336424 326262
rect 336372 326198 336424 326204
rect 335648 321526 335860 321554
rect 335544 4956 335596 4962
rect 335544 4898 335596 4904
rect 335648 4894 335676 321526
rect 337580 316034 337608 338014
rect 338132 335782 338160 338014
rect 338120 335776 338172 335782
rect 338120 335718 338172 335724
rect 338212 326392 338264 326398
rect 338212 326334 338264 326340
rect 336936 316006 337608 316034
rect 336936 5030 336964 316006
rect 338224 5098 338252 326334
rect 338408 316034 338436 338014
rect 338776 326398 338804 338014
rect 339144 335646 339172 338014
rect 339604 336734 339632 338014
rect 339592 336728 339644 336734
rect 339592 336670 339644 336676
rect 339132 335640 339184 335646
rect 339132 335582 339184 335588
rect 338764 326392 338816 326398
rect 338764 326334 338816 326340
rect 339972 316034 340000 338014
rect 340432 335986 340460 338014
rect 340420 335980 340472 335986
rect 340420 335922 340472 335928
rect 338316 316006 338436 316034
rect 339604 316006 340000 316034
rect 338212 5092 338264 5098
rect 338212 5034 338264 5040
rect 336924 5024 336976 5030
rect 336924 4966 336976 4972
rect 335636 4888 335688 4894
rect 335636 4830 335688 4836
rect 336280 3936 336332 3942
rect 336280 3878 336332 3884
rect 335452 3868 335504 3874
rect 335452 3810 335504 3816
rect 333244 3460 333296 3466
rect 333244 3402 333296 3408
rect 333888 3460 333940 3466
rect 333888 3402 333940 3408
rect 334624 3460 334676 3466
rect 334624 3402 334676 3408
rect 333900 480 333928 3402
rect 335084 3324 335136 3330
rect 335084 3266 335136 3272
rect 335096 480 335124 3266
rect 336292 480 336320 3878
rect 337476 3868 337528 3874
rect 337476 3810 337528 3816
rect 337488 480 337516 3810
rect 338316 3126 338344 316006
rect 339604 5166 339632 316006
rect 339592 5160 339644 5166
rect 339592 5102 339644 5108
rect 340892 4298 340920 338014
rect 340972 330540 341024 330546
rect 340972 330482 341024 330488
rect 340800 4270 340920 4298
rect 340800 4078 340828 4270
rect 340984 4162 341012 330482
rect 341168 316034 341196 338014
rect 341628 330546 341656 338014
rect 342272 335918 342300 338014
rect 342260 335912 342312 335918
rect 342260 335854 342312 335860
rect 342456 335354 342484 338014
rect 342364 335326 342484 335354
rect 341616 330540 341668 330546
rect 341616 330482 341668 330488
rect 341076 316006 341196 316034
rect 341076 5234 341104 316006
rect 342364 5302 342392 335326
rect 342824 316034 342852 338014
rect 343192 336394 343220 338014
rect 343180 336388 343232 336394
rect 343180 336330 343232 336336
rect 342456 316006 342852 316034
rect 342352 5296 342404 5302
rect 342352 5238 342404 5244
rect 341064 5228 341116 5234
rect 341064 5170 341116 5176
rect 340892 4146 341012 4162
rect 340880 4140 341012 4146
rect 340932 4134 341012 4140
rect 342168 4140 342220 4146
rect 340880 4082 340932 4088
rect 342168 4082 342220 4088
rect 340788 4072 340840 4078
rect 340788 4014 340840 4020
rect 340972 4072 341024 4078
rect 340972 4014 341024 4020
rect 338672 4004 338724 4010
rect 338672 3946 338724 3952
rect 338304 3120 338356 3126
rect 338304 3062 338356 3068
rect 338684 480 338712 3946
rect 339868 3256 339920 3262
rect 339868 3198 339920 3204
rect 339880 480 339908 3198
rect 340984 480 341012 4014
rect 342180 480 342208 4082
rect 342456 3398 342484 316006
rect 343744 5370 343772 338014
rect 344020 316034 344048 338014
rect 344480 335850 344508 338014
rect 345032 336462 345060 338014
rect 345308 336818 345336 338014
rect 345124 336790 345336 336818
rect 345020 336456 345072 336462
rect 345020 336398 345072 336404
rect 344468 335844 344520 335850
rect 344468 335786 344520 335792
rect 343836 316006 344048 316034
rect 343732 5364 343784 5370
rect 343732 5306 343784 5312
rect 342444 3392 342496 3398
rect 342444 3334 342496 3340
rect 343364 3188 343416 3194
rect 343364 3130 343416 3136
rect 343376 480 343404 3130
rect 343836 3058 343864 316006
rect 345124 3534 345152 336790
rect 345676 336682 345704 338014
rect 345216 336654 345704 336682
rect 345216 3602 345244 336654
rect 345388 336592 345440 336598
rect 345388 336534 345440 336540
rect 345296 330540 345348 330546
rect 345296 330482 345348 330488
rect 345308 5438 345336 330482
rect 345296 5432 345348 5438
rect 345296 5374 345348 5380
rect 345204 3596 345256 3602
rect 345204 3538 345256 3544
rect 345112 3528 345164 3534
rect 345112 3470 345164 3476
rect 344560 3460 344612 3466
rect 344560 3402 344612 3408
rect 343824 3052 343876 3058
rect 343824 2994 343876 3000
rect 344572 480 344600 3402
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345400 354 345428 336534
rect 346044 330546 346072 338014
rect 346032 330540 346084 330546
rect 346032 330482 346084 330488
rect 346504 3670 346532 338014
rect 346872 336190 346900 338014
rect 347332 336326 347360 338014
rect 347320 336320 347372 336326
rect 347320 336262 347372 336268
rect 347792 336258 347820 338014
rect 347780 336252 347832 336258
rect 347780 336194 347832 336200
rect 346860 336184 346912 336190
rect 346860 336126 346912 336132
rect 348068 316034 348096 338014
rect 348528 336054 348556 338014
rect 348516 336048 348568 336054
rect 348516 335990 348568 335996
rect 349448 335354 349476 338014
rect 349540 338014 349600 338042
rect 349724 338014 349968 338042
rect 350092 338014 350428 338042
rect 350644 338014 350796 338042
rect 350920 338014 351256 338042
rect 351380 338014 351624 338042
rect 352084 338014 352236 338042
rect 349540 336122 349568 338014
rect 349528 336116 349580 336122
rect 349528 336058 349580 336064
rect 349448 335326 349568 335354
rect 349344 330540 349396 330546
rect 349344 330482 349396 330488
rect 349252 330268 349304 330274
rect 349252 330210 349304 330216
rect 347884 316006 348096 316034
rect 347884 3738 347912 316006
rect 349264 3942 349292 330210
rect 349252 3936 349304 3942
rect 349252 3878 349304 3884
rect 347872 3732 347924 3738
rect 347872 3674 347924 3680
rect 346492 3664 346544 3670
rect 346492 3606 346544 3612
rect 349252 3664 349304 3670
rect 349252 3606 349304 3612
rect 348056 3392 348108 3398
rect 348056 3334 348108 3340
rect 346952 3324 347004 3330
rect 346952 3266 347004 3272
rect 346964 480 346992 3266
rect 348068 480 348096 3334
rect 349264 480 349292 3606
rect 349356 3466 349384 330482
rect 349540 3806 349568 335326
rect 349724 330546 349752 338014
rect 349712 330540 349764 330546
rect 349712 330482 349764 330488
rect 350092 330274 350120 338014
rect 350080 330268 350132 330274
rect 350080 330210 350132 330216
rect 350540 326392 350592 326398
rect 350540 326334 350592 326340
rect 349528 3800 349580 3806
rect 349528 3742 349580 3748
rect 349344 3460 349396 3466
rect 349344 3402 349396 3408
rect 350552 3262 350580 326334
rect 350644 3874 350672 338014
rect 350920 316034 350948 338014
rect 351380 326398 351408 338014
rect 352208 328454 352236 338014
rect 352116 328426 352236 328454
rect 352300 338014 352452 338042
rect 352576 338014 352820 338042
rect 352944 338014 353280 338042
rect 353404 338014 353648 338042
rect 353772 338014 354108 338042
rect 354232 338014 354476 338042
rect 352012 326460 352064 326466
rect 352012 326402 352064 326408
rect 351368 326392 351420 326398
rect 351368 326334 351420 326340
rect 351920 326392 351972 326398
rect 351920 326334 351972 326340
rect 350736 316006 350948 316034
rect 350736 4010 350764 316006
rect 351644 4072 351696 4078
rect 351644 4014 351696 4020
rect 350724 4004 350776 4010
rect 350724 3946 350776 3952
rect 350632 3868 350684 3874
rect 350632 3810 350684 3816
rect 350540 3256 350592 3262
rect 350540 3198 350592 3204
rect 350448 3052 350500 3058
rect 350448 2994 350500 3000
rect 350460 480 350488 2994
rect 351656 480 351684 4014
rect 351932 3194 351960 326334
rect 352024 3534 352052 326402
rect 352116 323762 352144 328426
rect 352116 323734 352236 323762
rect 352104 323604 352156 323610
rect 352104 323546 352156 323552
rect 352116 4146 352144 323546
rect 352104 4140 352156 4146
rect 352104 4082 352156 4088
rect 352208 4010 352236 323734
rect 352300 323610 352328 338014
rect 352576 326398 352604 338014
rect 352944 326466 352972 338014
rect 353404 336598 353432 338014
rect 353392 336592 353444 336598
rect 353392 336534 353444 336540
rect 353772 335354 353800 338014
rect 353404 335326 353800 335354
rect 353944 335368 353996 335374
rect 352932 326460 352984 326466
rect 352932 326402 352984 326408
rect 352564 326392 352616 326398
rect 352564 326334 352616 326340
rect 352288 323604 352340 323610
rect 352288 323546 352340 323552
rect 352196 4004 352248 4010
rect 352196 3946 352248 3952
rect 352012 3528 352064 3534
rect 352012 3470 352064 3476
rect 352840 3528 352892 3534
rect 352840 3470 352892 3476
rect 351920 3188 351972 3194
rect 351920 3130 351972 3136
rect 352852 480 352880 3470
rect 353404 3330 353432 335326
rect 353944 335310 353996 335316
rect 353484 326392 353536 326398
rect 353484 326334 353536 326340
rect 353496 3398 353524 326334
rect 353956 3534 353984 335310
rect 354232 326398 354260 338014
rect 354830 337770 354858 338028
rect 354968 338014 355304 338042
rect 355428 338014 355672 338042
rect 356072 338014 356132 338042
rect 356256 338014 356500 338042
rect 356624 338014 356868 338042
rect 356992 338014 357328 338042
rect 357452 338014 357696 338042
rect 357820 338014 358156 338042
rect 358524 338014 358768 338042
rect 354830 337742 354904 337770
rect 354680 336728 354732 336734
rect 354680 336670 354732 336676
rect 354220 326392 354272 326398
rect 354220 326334 354272 326340
rect 353944 3528 353996 3534
rect 353944 3470 353996 3476
rect 353484 3392 353536 3398
rect 353484 3334 353536 3340
rect 353392 3324 353444 3330
rect 353392 3266 353444 3272
rect 354036 3324 354088 3330
rect 354036 3266 354088 3272
rect 354048 480 354076 3266
rect 354692 3058 354720 336670
rect 354772 326392 354824 326398
rect 354772 326334 354824 326340
rect 354784 4078 354812 326334
rect 354772 4072 354824 4078
rect 354772 4014 354824 4020
rect 354876 3670 354904 337742
rect 354968 336734 354996 338014
rect 354956 336728 355008 336734
rect 354956 336670 355008 336676
rect 355428 326398 355456 338014
rect 356072 335374 356100 338014
rect 356256 336682 356284 338014
rect 356164 336654 356284 336682
rect 356060 335368 356112 335374
rect 356060 335310 356112 335316
rect 355416 326392 355468 326398
rect 355416 326334 355468 326340
rect 354864 3664 354916 3670
rect 354864 3606 354916 3612
rect 355232 3528 355284 3534
rect 355232 3470 355284 3476
rect 354680 3052 354732 3058
rect 354680 2994 354732 3000
rect 355244 480 355272 3470
rect 356164 3330 356192 336654
rect 356624 335354 356652 338014
rect 356256 335326 356652 335354
rect 356256 3534 356284 335326
rect 356992 316034 357020 338014
rect 356348 316006 357020 316034
rect 356244 3528 356296 3534
rect 356244 3470 356296 3476
rect 356152 3324 356204 3330
rect 356152 3266 356204 3272
rect 356348 480 356376 316006
rect 357452 3346 357480 338014
rect 357820 316034 357848 338014
rect 358740 335354 358768 338014
rect 358878 337770 358906 338028
rect 359016 338014 359352 338042
rect 359720 338014 360056 338042
rect 358878 337742 358952 337770
rect 358740 335326 358860 335354
rect 357544 316006 357848 316034
rect 357544 3534 357572 316006
rect 357532 3528 357584 3534
rect 357532 3470 357584 3476
rect 358728 3528 358780 3534
rect 358728 3470 358780 3476
rect 357452 3318 357572 3346
rect 357544 480 357572 3318
rect 358740 480 358768 3470
rect 358832 626 358860 335326
rect 358924 3534 358952 337742
rect 358912 3528 358964 3534
rect 358912 3470 358964 3476
rect 359016 3194 359044 338014
rect 360028 336666 360056 338014
rect 360120 338014 360180 338042
rect 360396 338014 360548 338042
rect 360672 338014 361008 338042
rect 361132 338014 361376 338042
rect 361592 338014 361744 338042
rect 362144 338014 362204 338042
rect 362328 338014 362572 338042
rect 360120 336734 360148 338014
rect 360108 336728 360160 336734
rect 360108 336670 360160 336676
rect 360016 336660 360068 336666
rect 360016 336602 360068 336608
rect 360292 330540 360344 330546
rect 360292 330482 360344 330488
rect 360200 330472 360252 330478
rect 360200 330414 360252 330420
rect 360212 3738 360240 330414
rect 360304 4010 360332 330482
rect 360292 4004 360344 4010
rect 360292 3946 360344 3952
rect 360200 3732 360252 3738
rect 360200 3674 360252 3680
rect 359004 3188 359056 3194
rect 359004 3130 359056 3136
rect 360396 3058 360424 338014
rect 360672 330546 360700 338014
rect 360844 336728 360896 336734
rect 360844 336670 360896 336676
rect 360660 330540 360712 330546
rect 360660 330482 360712 330488
rect 360856 4078 360884 336670
rect 361132 330478 361160 338014
rect 361120 330472 361172 330478
rect 361120 330414 361172 330420
rect 360844 4072 360896 4078
rect 360844 4014 360896 4020
rect 361592 3670 361620 338014
rect 362144 335850 362172 338014
rect 362132 335844 362184 335850
rect 362132 335786 362184 335792
rect 362328 316034 362356 338014
rect 363018 337770 363046 338028
rect 363156 338014 363400 338042
rect 363524 338014 363768 338042
rect 363892 338014 364228 338042
rect 364352 338014 364596 338042
rect 364996 338014 365056 338042
rect 365180 338014 365424 338042
rect 363018 337742 363092 337770
rect 362960 336660 363012 336666
rect 362960 336602 363012 336608
rect 361684 316006 362356 316034
rect 361580 3664 361632 3670
rect 361580 3606 361632 3612
rect 361120 3528 361172 3534
rect 361120 3470 361172 3476
rect 360384 3052 360436 3058
rect 360384 2994 360436 3000
rect 358832 598 359504 626
rect 345726 354 345838 480
rect 345400 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 598
rect 361132 480 361160 3470
rect 361684 3398 361712 316006
rect 362972 3482 363000 336602
rect 363064 330546 363092 337742
rect 363052 330540 363104 330546
rect 363052 330482 363104 330488
rect 363052 328364 363104 328370
rect 363052 328306 363104 328312
rect 363064 3874 363092 328306
rect 363156 3942 363184 338014
rect 363524 335354 363552 338014
rect 363604 335844 363656 335850
rect 363604 335786 363656 335792
rect 363248 335326 363552 335354
rect 363248 4146 363276 335326
rect 363328 330540 363380 330546
rect 363328 330482 363380 330488
rect 363236 4140 363288 4146
rect 363236 4082 363288 4088
rect 363144 3936 363196 3942
rect 363144 3878 363196 3884
rect 363052 3868 363104 3874
rect 363052 3810 363104 3816
rect 363340 3806 363368 330482
rect 363328 3800 363380 3806
rect 363328 3742 363380 3748
rect 362972 3454 363552 3482
rect 361672 3392 361724 3398
rect 361672 3334 361724 3340
rect 362316 3188 362368 3194
rect 362316 3130 362368 3136
rect 362328 480 362356 3130
rect 363524 480 363552 3454
rect 363616 3194 363644 335786
rect 363892 328370 363920 338014
rect 363880 328364 363932 328370
rect 363880 328306 363932 328312
rect 363696 3800 363748 3806
rect 363696 3742 363748 3748
rect 363708 3262 363736 3742
rect 364352 3534 364380 338014
rect 364996 336598 365024 338014
rect 364984 336592 365036 336598
rect 364984 336534 365036 336540
rect 365180 316034 365208 338014
rect 365778 337770 365806 338028
rect 366252 338014 366496 338042
rect 366620 338014 366864 338042
rect 365778 337742 365852 337770
rect 365720 328772 365772 328778
rect 365720 328714 365772 328720
rect 364444 316006 365208 316034
rect 364340 3528 364392 3534
rect 364340 3470 364392 3476
rect 364444 3466 364472 316006
rect 365732 4078 365760 328714
rect 364616 4072 364668 4078
rect 364616 4014 364668 4020
rect 365720 4072 365772 4078
rect 365720 4014 365772 4020
rect 364432 3460 364484 3466
rect 364432 3402 364484 3408
rect 363696 3256 363748 3262
rect 363696 3198 363748 3204
rect 363604 3188 363656 3194
rect 363604 3130 363656 3136
rect 364628 480 364656 4014
rect 365824 3738 365852 337742
rect 366468 336530 366496 338014
rect 366456 336524 366508 336530
rect 366456 336466 366508 336472
rect 366836 336054 366864 338014
rect 366928 338014 367080 338042
rect 367204 338014 367448 338042
rect 367572 338014 367816 338042
rect 367940 338014 368276 338042
rect 368584 338014 368644 338042
rect 368768 338014 369104 338042
rect 369472 338014 369808 338042
rect 366824 336048 366876 336054
rect 366824 335990 366876 335996
rect 366928 328778 366956 338014
rect 367204 335354 367232 338014
rect 367112 335326 367232 335354
rect 366916 328772 366968 328778
rect 366916 328714 366968 328720
rect 367112 5098 367140 335326
rect 367192 330540 367244 330546
rect 367192 330482 367244 330488
rect 367100 5092 367152 5098
rect 367100 5034 367152 5040
rect 367204 4146 367232 330482
rect 367572 316034 367600 338014
rect 367940 330546 367968 338014
rect 368584 336394 368612 338014
rect 368572 336388 368624 336394
rect 368572 336330 368624 336336
rect 367928 330540 367980 330546
rect 367928 330482 367980 330488
rect 368768 316034 368796 338014
rect 369780 336734 369808 338014
rect 369872 338014 369932 338042
rect 370056 338014 370300 338042
rect 370668 338014 371004 338042
rect 369768 336728 369820 336734
rect 369768 336670 369820 336676
rect 369872 336326 369900 338014
rect 369860 336320 369912 336326
rect 369860 336262 369912 336268
rect 370056 316034 370084 338014
rect 370976 335918 371004 338014
rect 371068 338014 371128 338042
rect 371252 338014 371496 338042
rect 371896 338014 371956 338042
rect 372080 338014 372324 338042
rect 372692 338014 373028 338042
rect 373152 338014 373396 338042
rect 373520 338014 373764 338042
rect 371068 336258 371096 338014
rect 371056 336252 371108 336258
rect 371056 336194 371108 336200
rect 370964 335912 371016 335918
rect 370964 335854 371016 335860
rect 367296 316006 367600 316034
rect 368492 316006 368796 316034
rect 369872 316006 370084 316034
rect 367296 5234 367324 316006
rect 367284 5228 367336 5234
rect 367284 5170 367336 5176
rect 367284 5092 367336 5098
rect 367284 5034 367336 5040
rect 367100 4140 367152 4146
rect 367100 4082 367152 4088
rect 367192 4140 367244 4146
rect 367192 4082 367244 4088
rect 367008 4004 367060 4010
rect 367008 3946 367060 3952
rect 365812 3732 365864 3738
rect 365812 3674 365864 3680
rect 365812 3052 365864 3058
rect 365812 2994 365864 3000
rect 365824 480 365852 2994
rect 367020 480 367048 3946
rect 367112 3806 367140 4082
rect 367100 3800 367152 3806
rect 367100 3742 367152 3748
rect 367296 3330 367324 5034
rect 368492 4010 368520 316006
rect 368480 4004 368532 4010
rect 368480 3946 368532 3952
rect 368204 3664 368256 3670
rect 368204 3606 368256 3612
rect 367284 3324 367336 3330
rect 367284 3266 367336 3272
rect 368216 480 368244 3606
rect 369400 3596 369452 3602
rect 369400 3538 369452 3544
rect 369412 480 369440 3538
rect 369872 3126 369900 316006
rect 370872 3868 370924 3874
rect 370872 3810 370924 3816
rect 370884 3670 370912 3810
rect 370872 3664 370924 3670
rect 370872 3606 370924 3612
rect 371252 3602 371280 338014
rect 371896 335442 371924 338014
rect 371884 335436 371936 335442
rect 371884 335378 371936 335384
rect 372080 316034 372108 338014
rect 373000 336190 373028 338014
rect 373368 336734 373396 338014
rect 373264 336728 373316 336734
rect 373264 336670 373316 336676
rect 373356 336728 373408 336734
rect 373356 336670 373408 336676
rect 372988 336184 373040 336190
rect 372988 336126 373040 336132
rect 371344 316006 372108 316034
rect 371344 5166 371372 316006
rect 371332 5160 371384 5166
rect 371332 5102 371384 5108
rect 371240 3596 371292 3602
rect 371240 3538 371292 3544
rect 371700 3392 371752 3398
rect 371700 3334 371752 3340
rect 370596 3188 370648 3194
rect 370596 3130 370648 3136
rect 369860 3120 369912 3126
rect 369860 3062 369912 3068
rect 370608 480 370636 3130
rect 371712 480 371740 3334
rect 372896 3256 372948 3262
rect 372896 3198 372948 3204
rect 372908 480 372936 3198
rect 373276 3058 373304 336670
rect 373736 336666 373764 338014
rect 373920 338014 373980 338042
rect 374288 338014 374348 338042
rect 374472 338014 374716 338042
rect 375176 338014 375328 338042
rect 373724 336660 373776 336666
rect 373724 336602 373776 336608
rect 373920 335986 373948 338014
rect 373908 335980 373960 335986
rect 373908 335922 373960 335928
rect 374288 335714 374316 338014
rect 374276 335708 374328 335714
rect 374276 335650 374328 335656
rect 374472 316034 374500 338014
rect 375300 336462 375328 338014
rect 375484 338014 375544 338042
rect 375668 338014 376004 338042
rect 376372 338014 376616 338042
rect 375288 336456 375340 336462
rect 375288 336398 375340 336404
rect 374736 336048 374788 336054
rect 374736 335990 374788 335996
rect 374644 335912 374696 335918
rect 374644 335854 374696 335860
rect 374012 316006 374500 316034
rect 374012 5098 374040 316006
rect 374000 5092 374052 5098
rect 374000 5034 374052 5040
rect 374092 3868 374144 3874
rect 374092 3810 374144 3816
rect 373264 3052 373316 3058
rect 373264 2994 373316 3000
rect 374104 480 374132 3810
rect 374656 3194 374684 335854
rect 374748 3262 374776 335990
rect 375484 335782 375512 338014
rect 375472 335776 375524 335782
rect 375472 335718 375524 335724
rect 375668 316034 375696 338014
rect 376588 336054 376616 338014
rect 376680 338014 376740 338042
rect 376864 338014 377200 338042
rect 377568 338014 377904 338042
rect 376576 336048 376628 336054
rect 376576 335990 376628 335996
rect 376680 335850 376708 338014
rect 376668 335844 376720 335850
rect 376668 335786 376720 335792
rect 376024 335436 376076 335442
rect 376024 335378 376076 335384
rect 375392 316006 375696 316034
rect 375392 5030 375420 316006
rect 375380 5024 375432 5030
rect 375380 4966 375432 4972
rect 376036 3806 376064 335378
rect 376864 316034 376892 338014
rect 377404 336592 377456 336598
rect 377404 336534 377456 336540
rect 376772 316006 376892 316034
rect 376772 4962 376800 316006
rect 376760 4956 376812 4962
rect 376760 4898 376812 4904
rect 377416 4010 377444 336534
rect 377876 336025 377904 338014
rect 377968 338014 378028 338042
rect 378244 338014 378396 338042
rect 378520 338014 378856 338042
rect 378980 338014 379224 338042
rect 379532 338014 379592 338042
rect 377968 336122 377996 338014
rect 378140 336728 378192 336734
rect 378140 336670 378192 336676
rect 377956 336116 378008 336122
rect 377956 336058 378008 336064
rect 377862 336016 377918 336025
rect 377862 335951 377918 335960
rect 378152 4486 378180 336670
rect 378244 4894 378272 338014
rect 378520 336734 378548 338014
rect 378508 336728 378560 336734
rect 378508 336670 378560 336676
rect 378980 316034 379008 338014
rect 378336 316006 379008 316034
rect 378232 4888 378284 4894
rect 378232 4830 378284 4836
rect 378336 4826 378364 316006
rect 378324 4820 378376 4826
rect 378324 4762 378376 4768
rect 379532 4554 379560 338014
rect 380038 337770 380066 338028
rect 380176 338014 380420 338042
rect 380544 338014 380880 338042
rect 381004 338014 381248 338042
rect 381372 338014 381616 338042
rect 381740 338014 382076 338042
rect 382384 338014 382444 338042
rect 382568 338014 382904 338042
rect 383028 338014 383272 338042
rect 383396 338014 383640 338042
rect 383764 338014 384100 338042
rect 384224 338014 384468 338042
rect 384592 338014 384928 338042
rect 385052 338014 385296 338042
rect 385420 338014 385756 338042
rect 386124 338014 386368 338042
rect 386492 338014 386644 338042
rect 380038 337742 380112 337770
rect 379980 336524 380032 336530
rect 379980 336466 380032 336472
rect 379992 335354 380020 336466
rect 380084 335986 380112 337742
rect 380072 335980 380124 335986
rect 380072 335922 380124 335928
rect 379992 335326 380112 335354
rect 379612 330540 379664 330546
rect 379612 330482 379664 330488
rect 379624 4622 379652 330482
rect 379704 330472 379756 330478
rect 379704 330414 379756 330420
rect 379716 6390 379744 330414
rect 380084 325694 380112 335326
rect 380176 330546 380204 338014
rect 380256 336728 380308 336734
rect 380256 336670 380308 336676
rect 380164 330540 380216 330546
rect 380164 330482 380216 330488
rect 380084 325666 380204 325694
rect 379704 6384 379756 6390
rect 379704 6326 379756 6332
rect 379612 4616 379664 4622
rect 379612 4558 379664 4564
rect 379520 4548 379572 4554
rect 379520 4490 379572 4496
rect 378140 4480 378192 4486
rect 378140 4422 378192 4428
rect 378796 4146 379008 4162
rect 378784 4140 379008 4146
rect 378836 4134 379008 4140
rect 378784 4082 378836 4088
rect 378980 4010 379008 4134
rect 377404 4004 377456 4010
rect 377404 3946 377456 3952
rect 378876 4004 378928 4010
rect 378876 3946 378928 3952
rect 378968 4004 379020 4010
rect 378968 3946 379020 3952
rect 375288 3800 375340 3806
rect 375288 3742 375340 3748
rect 376024 3800 376076 3806
rect 376024 3742 376076 3748
rect 374736 3256 374788 3262
rect 374736 3198 374788 3204
rect 374644 3188 374696 3194
rect 374644 3130 374696 3136
rect 375300 480 375328 3742
rect 376484 3664 376536 3670
rect 376484 3606 376536 3612
rect 376576 3664 376628 3670
rect 376576 3606 376628 3612
rect 376496 480 376524 3606
rect 376588 3126 376616 3606
rect 377680 3528 377732 3534
rect 377680 3470 377732 3476
rect 376576 3120 376628 3126
rect 376576 3062 376628 3068
rect 377692 480 377720 3470
rect 378888 480 378916 3946
rect 379980 3392 380032 3398
rect 379980 3334 380032 3340
rect 380072 3392 380124 3398
rect 380072 3334 380124 3340
rect 379992 480 380020 3334
rect 380084 3194 380112 3334
rect 380072 3188 380124 3194
rect 380072 3130 380124 3136
rect 380176 2990 380204 325666
rect 380268 3534 380296 336670
rect 380544 330478 380572 338014
rect 381004 336682 381032 338014
rect 380912 336654 381032 336682
rect 380532 330472 380584 330478
rect 380532 330414 380584 330420
rect 380256 3528 380308 3534
rect 380256 3470 380308 3476
rect 380912 3194 380940 336654
rect 381372 335354 381400 338014
rect 381004 335326 381400 335354
rect 381004 6322 381032 335326
rect 381740 316034 381768 338014
rect 382280 330472 382332 330478
rect 382280 330414 382332 330420
rect 381096 316006 381768 316034
rect 380992 6316 381044 6322
rect 380992 6258 381044 6264
rect 381096 6254 381124 316006
rect 381084 6248 381136 6254
rect 381084 6190 381136 6196
rect 382292 3942 382320 330414
rect 382280 3936 382332 3942
rect 382280 3878 382332 3884
rect 381176 3732 381228 3738
rect 381176 3674 381228 3680
rect 380900 3188 380952 3194
rect 380900 3130 380952 3136
rect 380164 2984 380216 2990
rect 380164 2926 380216 2932
rect 381188 480 381216 3674
rect 382384 3466 382412 338014
rect 382464 330540 382516 330546
rect 382464 330482 382516 330488
rect 382476 5846 382504 330482
rect 382568 5914 382596 338014
rect 383028 330546 383056 338014
rect 383016 330540 383068 330546
rect 383016 330482 383068 330488
rect 383396 330478 383424 338014
rect 383660 330540 383712 330546
rect 383660 330482 383712 330488
rect 383384 330472 383436 330478
rect 383384 330414 383436 330420
rect 382556 5908 382608 5914
rect 382556 5850 382608 5856
rect 382464 5840 382516 5846
rect 382464 5782 382516 5788
rect 383672 4146 383700 330482
rect 383764 6526 383792 338014
rect 384224 316034 384252 338014
rect 384304 336388 384356 336394
rect 384304 336330 384356 336336
rect 383856 316006 384252 316034
rect 383856 8770 383884 316006
rect 383844 8764 383896 8770
rect 383844 8706 383896 8712
rect 383752 6520 383804 6526
rect 383752 6462 383804 6468
rect 383660 4140 383712 4146
rect 383660 4082 383712 4088
rect 382372 3460 382424 3466
rect 382372 3402 382424 3408
rect 384316 3262 384344 336330
rect 384592 330546 384620 338014
rect 384580 330540 384632 330546
rect 384580 330482 384632 330488
rect 385052 5982 385080 338014
rect 385420 316034 385448 338014
rect 386340 336734 386368 338014
rect 386328 336728 386380 336734
rect 386328 336670 386380 336676
rect 386512 330540 386564 330546
rect 386512 330482 386564 330488
rect 385144 316006 385448 316034
rect 385144 8838 385172 316006
rect 385132 8832 385184 8838
rect 385132 8774 385184 8780
rect 386524 6118 386552 330482
rect 386512 6112 386564 6118
rect 386512 6054 386564 6060
rect 386616 6050 386644 338014
rect 386708 338014 386952 338042
rect 387076 338014 387320 338042
rect 387444 338014 387780 338042
rect 387904 338014 388148 338042
rect 388456 338014 388516 338042
rect 388640 338014 388976 338042
rect 389284 338014 389344 338042
rect 389744 338014 389804 338042
rect 389928 338014 390172 338042
rect 390296 338014 390540 338042
rect 390756 338014 391000 338042
rect 391124 338014 391368 338042
rect 391492 338014 391828 338042
rect 391952 338014 392196 338042
rect 392320 338014 392564 338042
rect 392688 338014 393024 338042
rect 393332 338014 393392 338042
rect 393516 338014 393852 338042
rect 393976 338014 394220 338042
rect 394620 338014 394680 338042
rect 394804 338014 395048 338042
rect 395172 338014 395416 338042
rect 395876 338014 396028 338042
rect 396244 338014 396396 338042
rect 386708 8906 386736 338014
rect 387076 335354 387104 338014
rect 387156 335708 387208 335714
rect 387156 335650 387208 335656
rect 386984 335326 387104 335354
rect 386984 316034 387012 335326
rect 387168 316034 387196 335650
rect 387444 330546 387472 338014
rect 387432 330540 387484 330546
rect 387432 330482 387484 330488
rect 387800 329588 387852 329594
rect 387800 329530 387852 329536
rect 386800 316006 387012 316034
rect 387076 316006 387196 316034
rect 386696 8900 386748 8906
rect 386696 8842 386748 8848
rect 386604 6044 386656 6050
rect 386604 5986 386656 5992
rect 385040 5976 385092 5982
rect 385040 5918 385092 5924
rect 384764 4072 384816 4078
rect 384764 4014 384816 4020
rect 383568 3256 383620 3262
rect 383568 3198 383620 3204
rect 384304 3256 384356 3262
rect 384304 3198 384356 3204
rect 382372 2984 382424 2990
rect 382372 2926 382424 2932
rect 382384 480 382412 2926
rect 383580 480 383608 3198
rect 384776 480 384804 4014
rect 386800 3369 386828 316006
rect 386786 3360 386842 3369
rect 385960 3324 386012 3330
rect 387076 3330 387104 316006
rect 387812 6866 387840 329530
rect 387904 9654 387932 338014
rect 388456 336598 388484 338014
rect 388444 336592 388496 336598
rect 388444 336534 388496 336540
rect 388444 336320 388496 336326
rect 388444 336262 388496 336268
rect 387892 9648 387944 9654
rect 387892 9590 387944 9596
rect 387800 6860 387852 6866
rect 387800 6802 387852 6808
rect 387156 5228 387208 5234
rect 387156 5170 387208 5176
rect 386786 3295 386842 3304
rect 387064 3324 387116 3330
rect 385960 3266 386012 3272
rect 387064 3266 387116 3272
rect 385972 480 386000 3266
rect 387168 480 387196 5170
rect 388352 4140 388404 4146
rect 388352 4082 388404 4088
rect 388260 4004 388312 4010
rect 388260 3946 388312 3952
rect 388272 480 388300 3946
rect 388364 3534 388392 4082
rect 388456 3738 388484 336262
rect 388640 329594 388668 338014
rect 388628 329588 388680 329594
rect 388628 329530 388680 329536
rect 389180 322516 389232 322522
rect 389180 322458 389232 322464
rect 389192 6798 389220 322458
rect 389284 9586 389312 338014
rect 389744 336530 389772 338014
rect 389732 336524 389784 336530
rect 389732 336466 389784 336472
rect 389824 335776 389876 335782
rect 389824 335718 389876 335724
rect 389364 326392 389416 326398
rect 389364 326334 389416 326340
rect 389272 9580 389324 9586
rect 389272 9522 389324 9528
rect 389376 9518 389404 326334
rect 389364 9512 389416 9518
rect 389364 9454 389416 9460
rect 389180 6792 389232 6798
rect 389180 6734 389232 6740
rect 388444 3732 388496 3738
rect 388444 3674 388496 3680
rect 388352 3528 388404 3534
rect 388352 3470 388404 3476
rect 388444 3528 388496 3534
rect 388444 3470 388496 3476
rect 388456 3194 388484 3470
rect 389456 3256 389508 3262
rect 389456 3198 389508 3204
rect 388444 3188 388496 3194
rect 388444 3130 388496 3136
rect 389468 480 389496 3198
rect 389836 3194 389864 335718
rect 389928 322522 389956 338014
rect 390296 326398 390324 338014
rect 390284 326392 390336 326398
rect 390284 326334 390336 326340
rect 390652 325372 390704 325378
rect 390652 325314 390704 325320
rect 390560 323060 390612 323066
rect 390560 323002 390612 323008
rect 389916 322516 389968 322522
rect 389916 322458 389968 322464
rect 390572 6730 390600 323002
rect 390664 10198 390692 325314
rect 390756 12986 390784 338014
rect 391124 323066 391152 338014
rect 391204 335844 391256 335850
rect 391204 335786 391256 335792
rect 391112 323060 391164 323066
rect 391112 323002 391164 323008
rect 390744 12980 390796 12986
rect 390744 12922 390796 12928
rect 390652 10192 390704 10198
rect 390652 10134 390704 10140
rect 390560 6724 390612 6730
rect 390560 6666 390612 6672
rect 391216 4078 391244 335786
rect 391492 325378 391520 338014
rect 391480 325372 391532 325378
rect 391480 325314 391532 325320
rect 391204 4072 391256 4078
rect 391204 4014 391256 4020
rect 391952 3874 391980 338014
rect 392320 335354 392348 338014
rect 392044 335326 392348 335354
rect 392044 6662 392072 335326
rect 392688 316034 392716 338014
rect 393332 336326 393360 338014
rect 393320 336320 393372 336326
rect 393320 336262 393372 336268
rect 393516 335354 393544 338014
rect 393976 336682 394004 338014
rect 392136 316006 392716 316034
rect 393332 335326 393544 335354
rect 393792 336654 394004 336682
rect 392136 10266 392164 316006
rect 392124 10260 392176 10266
rect 392124 10202 392176 10208
rect 392032 6656 392084 6662
rect 392032 6598 392084 6604
rect 393332 6594 393360 335326
rect 393792 316034 393820 336654
rect 394620 336394 394648 338014
rect 394608 336388 394660 336394
rect 394608 336330 394660 336336
rect 393964 336184 394016 336190
rect 393964 336126 394016 336132
rect 393424 316006 393820 316034
rect 393424 11014 393452 316006
rect 393976 16574 394004 336126
rect 394700 326392 394752 326398
rect 394700 326334 394752 326340
rect 393976 16546 394372 16574
rect 393412 11008 393464 11014
rect 393412 10950 393464 10956
rect 393320 6588 393372 6594
rect 393320 6530 393372 6536
rect 393136 4004 393188 4010
rect 393136 3946 393188 3952
rect 390652 3868 390704 3874
rect 390652 3810 390704 3816
rect 391940 3868 391992 3874
rect 391940 3810 391992 3816
rect 389824 3188 389876 3194
rect 389824 3130 389876 3136
rect 390664 480 390692 3810
rect 393148 3738 393176 3946
rect 393044 3732 393096 3738
rect 393044 3674 393096 3680
rect 393136 3732 393188 3738
rect 393136 3674 393188 3680
rect 391848 3120 391900 3126
rect 391848 3062 391900 3068
rect 391860 480 391888 3062
rect 393056 480 393084 3674
rect 394344 3670 394372 16546
rect 394712 10946 394740 326334
rect 394804 11558 394832 338014
rect 395172 326398 395200 338014
rect 396000 336190 396028 338014
rect 396080 336252 396132 336258
rect 396080 336194 396132 336200
rect 395988 336184 396040 336190
rect 395988 336126 396040 336132
rect 395160 326392 395212 326398
rect 395160 326334 395212 326340
rect 394792 11552 394844 11558
rect 394792 11494 394844 11500
rect 394700 10940 394752 10946
rect 394700 10882 394752 10888
rect 394240 3664 394292 3670
rect 394240 3606 394292 3612
rect 394332 3664 394384 3670
rect 394332 3606 394384 3612
rect 394252 480 394280 3606
rect 395344 3392 395396 3398
rect 395344 3334 395396 3340
rect 395356 480 395384 3334
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 336194
rect 396368 326534 396396 338014
rect 396460 338014 396704 338042
rect 396828 338014 397072 338042
rect 397196 338014 397440 338042
rect 397564 338014 397900 338042
rect 398024 338014 398268 338042
rect 398392 338014 398728 338042
rect 398944 338014 399096 338042
rect 399404 338014 399464 338042
rect 399588 338014 399924 338042
rect 396356 326528 396408 326534
rect 396356 326470 396408 326476
rect 396172 326392 396224 326398
rect 396172 326334 396224 326340
rect 396184 3398 396212 326334
rect 396460 323626 396488 338014
rect 396540 326528 396592 326534
rect 396540 326470 396592 326476
rect 396276 323598 396488 323626
rect 396276 10878 396304 323598
rect 396552 318794 396580 326470
rect 396828 326398 396856 338014
rect 396816 326392 396868 326398
rect 396816 326334 396868 326340
rect 396368 318766 396580 318794
rect 396368 11626 396396 318766
rect 397196 316034 397224 338014
rect 397460 326392 397512 326398
rect 397460 326334 397512 326340
rect 396460 316006 397224 316034
rect 396460 11694 396488 316006
rect 396448 11688 396500 11694
rect 396448 11630 396500 11636
rect 396356 11620 396408 11626
rect 396356 11562 396408 11568
rect 396264 10872 396316 10878
rect 396264 10814 396316 10820
rect 396172 3392 396224 3398
rect 396172 3334 396224 3340
rect 397472 3330 397500 326334
rect 397564 10810 397592 338014
rect 397644 326460 397696 326466
rect 397644 326402 397696 326408
rect 397656 12442 397684 326402
rect 398024 326398 398052 338014
rect 398104 335912 398156 335918
rect 398104 335854 398156 335860
rect 398012 326392 398064 326398
rect 398012 326334 398064 326340
rect 397644 12436 397696 12442
rect 397644 12378 397696 12384
rect 397552 10804 397604 10810
rect 397552 10746 397604 10752
rect 398116 3602 398144 335854
rect 398392 326466 398420 338014
rect 398380 326460 398432 326466
rect 398380 326402 398432 326408
rect 398840 326392 398892 326398
rect 398840 326334 398892 326340
rect 398852 10606 398880 326334
rect 398944 10742 398972 338014
rect 399404 336258 399432 338014
rect 399392 336252 399444 336258
rect 399392 336194 399444 336200
rect 399588 326398 399616 338014
rect 400278 337770 400306 338028
rect 400416 338014 400752 338042
rect 400876 338014 401120 338042
rect 401244 338014 401488 338042
rect 401704 338014 401948 338042
rect 402072 338014 402316 338042
rect 402440 338014 402776 338042
rect 400278 337742 400352 337770
rect 399576 326392 399628 326398
rect 399576 326334 399628 326340
rect 400220 326392 400272 326398
rect 400220 326334 400272 326340
rect 400324 326346 400352 337742
rect 400416 326482 400444 338014
rect 400772 336660 400824 336666
rect 400772 336602 400824 336608
rect 400416 326454 400628 326482
rect 398932 10736 398984 10742
rect 398932 10678 398984 10684
rect 398840 10600 398892 10606
rect 398840 10542 398892 10548
rect 400232 7410 400260 326334
rect 400324 326318 400536 326346
rect 400404 326256 400456 326262
rect 400404 326198 400456 326204
rect 400312 324284 400364 324290
rect 400312 324226 400364 324232
rect 400324 10538 400352 324226
rect 400416 10674 400444 326198
rect 400508 12374 400536 326318
rect 400600 326262 400628 326454
rect 400588 326256 400640 326262
rect 400588 326198 400640 326204
rect 400784 321554 400812 336602
rect 400876 324290 400904 338014
rect 401244 326398 401272 338014
rect 401232 326392 401284 326398
rect 401232 326334 401284 326340
rect 401600 325780 401652 325786
rect 401600 325722 401652 325728
rect 400864 324284 400916 324290
rect 400864 324226 400916 324232
rect 400784 321526 400904 321554
rect 400496 12368 400548 12374
rect 400496 12310 400548 12316
rect 400404 10668 400456 10674
rect 400404 10610 400456 10616
rect 400312 10532 400364 10538
rect 400312 10474 400364 10480
rect 400220 7404 400272 7410
rect 400220 7346 400272 7352
rect 400128 5160 400180 5166
rect 400128 5102 400180 5108
rect 398932 3800 398984 3806
rect 398932 3742 398984 3748
rect 397736 3596 397788 3602
rect 397736 3538 397788 3544
rect 398104 3596 398156 3602
rect 398104 3538 398156 3544
rect 397460 3324 397512 3330
rect 397460 3266 397512 3272
rect 397748 480 397776 3538
rect 398944 480 398972 3742
rect 400140 480 400168 5102
rect 400876 4214 400904 321526
rect 401612 7478 401640 325722
rect 401704 10470 401732 338014
rect 402072 316034 402100 338014
rect 402244 336456 402296 336462
rect 402244 336398 402296 336404
rect 401796 316006 402100 316034
rect 401692 10464 401744 10470
rect 401692 10406 401744 10412
rect 401796 10402 401824 316006
rect 402256 16574 402284 336398
rect 402440 325786 402468 338014
rect 403130 337770 403158 338028
rect 403268 338014 403604 338042
rect 403728 338014 403972 338042
rect 404096 338014 404340 338042
rect 404464 338014 404800 338042
rect 404924 338014 405168 338042
rect 405292 338014 405628 338042
rect 405752 338014 405996 338042
rect 406120 338014 406364 338042
rect 406488 338014 406824 338042
rect 407132 338014 407192 338042
rect 407316 338014 407652 338042
rect 407776 338014 408020 338042
rect 408144 338014 408388 338042
rect 408604 338014 408848 338042
rect 408972 338014 409216 338042
rect 409340 338014 409676 338042
rect 409984 338014 410044 338042
rect 410168 338014 410504 338042
rect 410628 338014 410872 338042
rect 410996 338014 411240 338042
rect 411456 338014 411700 338042
rect 411824 338014 412068 338042
rect 412192 338014 412528 338042
rect 412836 338014 412896 338042
rect 413020 338014 413264 338042
rect 413388 338014 413724 338042
rect 414092 338014 414336 338042
rect 403130 337742 403204 337770
rect 403176 328454 403204 337742
rect 403084 328426 403204 328454
rect 402980 326392 403032 326398
rect 402980 326334 403032 326340
rect 402428 325780 402480 325786
rect 402428 325722 402480 325728
rect 402256 16546 402652 16574
rect 401784 10396 401836 10402
rect 401784 10338 401836 10344
rect 401600 7472 401652 7478
rect 401600 7414 401652 7420
rect 400864 4208 400916 4214
rect 400864 4150 400916 4156
rect 402520 4140 402572 4146
rect 402520 4082 402572 4088
rect 401324 3664 401376 3670
rect 401324 3606 401376 3612
rect 401336 480 401364 3606
rect 402532 480 402560 4082
rect 402624 3806 402652 16546
rect 402992 7546 403020 326334
rect 403084 322810 403112 328426
rect 403084 322782 403204 322810
rect 403072 321700 403124 321706
rect 403072 321642 403124 321648
rect 403084 10334 403112 321642
rect 403176 12306 403204 322782
rect 403268 321706 403296 338014
rect 403728 326398 403756 338014
rect 403716 326392 403768 326398
rect 403716 326334 403768 326340
rect 403256 321700 403308 321706
rect 403256 321642 403308 321648
rect 404096 316034 404124 338014
rect 404360 326392 404412 326398
rect 404360 326334 404412 326340
rect 403268 316006 404124 316034
rect 403268 13054 403296 316006
rect 403256 13048 403308 13054
rect 403256 12990 403308 12996
rect 403164 12300 403216 12306
rect 403164 12242 403216 12248
rect 403072 10328 403124 10334
rect 403072 10270 403124 10276
rect 404372 8294 404400 326334
rect 404464 12238 404492 338014
rect 404544 326460 404596 326466
rect 404544 326402 404596 326408
rect 404556 13802 404584 326402
rect 404924 326398 404952 338014
rect 405004 336116 405056 336122
rect 405004 336058 405056 336064
rect 404912 326392 404964 326398
rect 404912 326334 404964 326340
rect 404544 13796 404596 13802
rect 404544 13738 404596 13744
rect 404452 12232 404504 12238
rect 404452 12174 404504 12180
rect 404360 8288 404412 8294
rect 404360 8230 404412 8236
rect 402980 7540 403032 7546
rect 402980 7482 403032 7488
rect 405016 4146 405044 336058
rect 405292 326466 405320 338014
rect 405280 326460 405332 326466
rect 405280 326402 405332 326408
rect 405752 4690 405780 338014
rect 406120 335354 406148 338014
rect 406384 335980 406436 335986
rect 406384 335922 406436 335928
rect 405844 335326 406148 335354
rect 405844 8226 405872 335326
rect 405924 326392 405976 326398
rect 405924 326334 405976 326340
rect 405936 13734 405964 326334
rect 405924 13728 405976 13734
rect 405924 13670 405976 13676
rect 405832 8220 405884 8226
rect 405832 8162 405884 8168
rect 405740 4684 405792 4690
rect 405740 4626 405792 4632
rect 403624 4140 403676 4146
rect 403624 4082 403676 4088
rect 405004 4140 405056 4146
rect 405004 4082 405056 4088
rect 402704 4004 402756 4010
rect 402704 3946 402756 3952
rect 402612 3800 402664 3806
rect 402612 3742 402664 3748
rect 402716 3602 402744 3946
rect 402704 3596 402756 3602
rect 402704 3538 402756 3544
rect 403636 480 403664 4082
rect 404820 4004 404872 4010
rect 404820 3946 404872 3952
rect 405740 4004 405792 4010
rect 405740 3946 405792 3952
rect 404832 480 404860 3946
rect 405752 3398 405780 3946
rect 406396 3670 406424 335922
rect 406488 326398 406516 338014
rect 406568 336048 406620 336054
rect 406568 335990 406620 335996
rect 406476 326392 406528 326398
rect 406476 326334 406528 326340
rect 406580 316034 406608 335990
rect 406488 316006 406608 316034
rect 406384 3664 406436 3670
rect 406384 3606 406436 3612
rect 406488 3602 406516 316006
rect 407132 4758 407160 338014
rect 407212 326392 407264 326398
rect 407212 326334 407264 326340
rect 407224 5506 407252 326334
rect 407316 8158 407344 338014
rect 407776 316034 407804 338014
rect 408144 326398 408172 338014
rect 408500 327344 408552 327350
rect 408500 327286 408552 327292
rect 408132 326392 408184 326398
rect 408132 326334 408184 326340
rect 407408 316006 407804 316034
rect 407408 13666 407436 316006
rect 407396 13660 407448 13666
rect 407396 13602 407448 13608
rect 407304 8152 407356 8158
rect 407304 8094 407356 8100
rect 407212 5500 407264 5506
rect 407212 5442 407264 5448
rect 408512 5438 408540 327286
rect 408604 8090 408632 338014
rect 408972 316034 409000 338014
rect 409142 336016 409198 336025
rect 409142 335951 409198 335960
rect 408696 316006 409000 316034
rect 408696 13598 408724 316006
rect 408684 13592 408736 13598
rect 408684 13534 408736 13540
rect 408592 8084 408644 8090
rect 408592 8026 408644 8032
rect 408500 5432 408552 5438
rect 408500 5374 408552 5380
rect 407212 5092 407264 5098
rect 407212 5034 407264 5040
rect 407120 4752 407172 4758
rect 407120 4694 407172 4700
rect 406476 3596 406528 3602
rect 406476 3538 406528 3544
rect 405740 3392 405792 3398
rect 405740 3334 405792 3340
rect 406016 3256 406068 3262
rect 406016 3198 406068 3204
rect 406028 480 406056 3198
rect 407224 480 407252 5034
rect 409156 3806 409184 335951
rect 409340 327350 409368 338014
rect 409880 330472 409932 330478
rect 409880 330414 409932 330420
rect 409328 327344 409380 327350
rect 409328 327286 409380 327292
rect 409892 5370 409920 330414
rect 409984 8022 410012 338014
rect 410064 330540 410116 330546
rect 410064 330482 410116 330488
rect 409972 8016 410024 8022
rect 409972 7958 410024 7964
rect 410076 7954 410104 330482
rect 410168 13530 410196 338014
rect 410628 330478 410656 338014
rect 410996 330546 411024 338014
rect 410984 330540 411036 330546
rect 410984 330482 411036 330488
rect 411260 330540 411312 330546
rect 411260 330482 411312 330488
rect 410616 330472 410668 330478
rect 410616 330414 410668 330420
rect 410156 13524 410208 13530
rect 410156 13466 410208 13472
rect 410064 7948 410116 7954
rect 410064 7890 410116 7896
rect 409880 5364 409932 5370
rect 409880 5306 409932 5312
rect 411272 5302 411300 330482
rect 411352 330472 411404 330478
rect 411352 330414 411404 330420
rect 411364 7886 411392 330414
rect 411456 13462 411484 338014
rect 411824 330546 411852 338014
rect 411904 336728 411956 336734
rect 411904 336670 411956 336676
rect 411812 330540 411864 330546
rect 411812 330482 411864 330488
rect 411916 16574 411944 336670
rect 412192 330478 412220 338014
rect 412836 335918 412864 338014
rect 412824 335912 412876 335918
rect 412824 335854 412876 335860
rect 413020 335354 413048 338014
rect 412652 335326 413048 335354
rect 412180 330472 412232 330478
rect 412180 330414 412232 330420
rect 411916 16546 412036 16574
rect 411444 13456 411496 13462
rect 411444 13398 411496 13404
rect 411352 7880 411404 7886
rect 411352 7822 411404 7828
rect 411260 5296 411312 5302
rect 411260 5238 411312 5244
rect 410800 5024 410852 5030
rect 410800 4966 410852 4972
rect 408408 3800 408460 3806
rect 408408 3742 408460 3748
rect 409144 3800 409196 3806
rect 409144 3742 409196 3748
rect 408420 480 408448 3742
rect 409604 3188 409656 3194
rect 409604 3130 409656 3136
rect 409616 480 409644 3130
rect 410812 480 410840 4966
rect 412008 4146 412036 16546
rect 412652 5234 412680 335326
rect 413388 316034 413416 338014
rect 414020 336728 414072 336734
rect 414020 336670 414072 336676
rect 412744 316006 413416 316034
rect 412744 7818 412772 316006
rect 412732 7812 412784 7818
rect 412732 7754 412784 7760
rect 412640 5228 412692 5234
rect 412640 5170 412692 5176
rect 414032 5166 414060 336670
rect 414112 330540 414164 330546
rect 414112 330482 414164 330488
rect 414124 7750 414152 330482
rect 414204 330472 414256 330478
rect 414204 330414 414256 330420
rect 414216 13326 414244 330414
rect 414308 13394 414336 338014
rect 414400 338014 414552 338042
rect 414676 338014 414920 338042
rect 415044 338014 415288 338042
rect 415412 338014 415748 338042
rect 415872 338014 416116 338042
rect 416576 338014 416728 338042
rect 414400 336734 414428 338014
rect 414388 336728 414440 336734
rect 414388 336670 414440 336676
rect 414676 330546 414704 338014
rect 414664 330540 414716 330546
rect 414664 330482 414716 330488
rect 415044 330478 415072 338014
rect 415032 330472 415084 330478
rect 415032 330414 415084 330420
rect 414296 13388 414348 13394
rect 414296 13330 414348 13336
rect 414204 13320 414256 13326
rect 414204 13262 414256 13268
rect 414112 7744 414164 7750
rect 414112 7686 414164 7692
rect 414020 5160 414072 5166
rect 414020 5102 414072 5108
rect 415412 5098 415440 338014
rect 415872 316034 415900 338014
rect 416044 336592 416096 336598
rect 416044 336534 416096 336540
rect 415504 316006 415900 316034
rect 415504 7682 415532 316006
rect 415492 7676 415544 7682
rect 415492 7618 415544 7624
rect 415400 5092 415452 5098
rect 415400 5034 415452 5040
rect 414296 4956 414348 4962
rect 414296 4898 414348 4904
rect 411904 4140 411956 4146
rect 411904 4082 411956 4088
rect 411996 4140 412048 4146
rect 411996 4082 412048 4088
rect 411916 3890 411944 4082
rect 413100 4072 413152 4078
rect 413100 4014 413152 4020
rect 411916 3862 412128 3890
rect 412100 3670 412128 3862
rect 412088 3664 412140 3670
rect 412088 3606 412140 3612
rect 411904 3596 411956 3602
rect 411904 3538 411956 3544
rect 411916 480 411944 3538
rect 413112 480 413140 4014
rect 414308 480 414336 4898
rect 416056 4078 416084 336534
rect 416700 336122 416728 338014
rect 416792 338014 416944 338042
rect 417068 338014 417312 338042
rect 417436 338014 417772 338042
rect 417896 338014 418140 338042
rect 418264 338014 418600 338042
rect 418908 338014 418968 338042
rect 419092 338014 419428 338042
rect 419736 338014 419796 338042
rect 419920 338014 420164 338042
rect 420288 338014 420624 338042
rect 416688 336116 416740 336122
rect 416688 336058 416740 336064
rect 416792 5030 416820 338014
rect 417068 335354 417096 338014
rect 416976 335326 417096 335354
rect 416872 329724 416924 329730
rect 416872 329666 416924 329672
rect 416780 5024 416832 5030
rect 416780 4966 416832 4972
rect 416884 4865 416912 329666
rect 416976 7614 417004 335326
rect 417436 316034 417464 338014
rect 417896 329730 417924 338014
rect 417884 329724 417936 329730
rect 417884 329666 417936 329672
rect 418160 326392 418212 326398
rect 418160 326334 418212 326340
rect 417068 316006 417464 316034
rect 417068 13258 417096 316006
rect 417056 13252 417108 13258
rect 417056 13194 417108 13200
rect 416964 7608 417016 7614
rect 416964 7550 417016 7556
rect 418172 4962 418200 326334
rect 418264 12170 418292 338014
rect 418908 336054 418936 338014
rect 418896 336048 418948 336054
rect 418896 335990 418948 335996
rect 419092 326398 419120 338014
rect 419736 326874 419764 338014
rect 419920 335354 419948 338014
rect 419828 335326 419948 335354
rect 419724 326868 419776 326874
rect 419724 326810 419776 326816
rect 419724 326664 419776 326670
rect 419724 326606 419776 326612
rect 419080 326392 419132 326398
rect 419080 326334 419132 326340
rect 419632 326392 419684 326398
rect 419632 326334 419684 326340
rect 419540 319252 419592 319258
rect 419540 319194 419592 319200
rect 418252 12164 418304 12170
rect 418252 12106 418304 12112
rect 418160 4956 418212 4962
rect 418160 4898 418212 4904
rect 417884 4888 417936 4894
rect 416870 4856 416926 4865
rect 417884 4830 417936 4836
rect 416870 4791 416926 4800
rect 416044 4072 416096 4078
rect 416044 4014 416096 4020
rect 415492 3800 415544 3806
rect 415492 3742 415544 3748
rect 415504 480 415532 3742
rect 416688 3664 416740 3670
rect 416688 3606 416740 3612
rect 416700 480 416728 3606
rect 417896 480 417924 4830
rect 418988 4480 419040 4486
rect 418988 4422 419040 4428
rect 419000 480 419028 4422
rect 419552 3806 419580 319194
rect 419644 4894 419672 326334
rect 419736 12102 419764 326606
rect 419828 319258 419856 335326
rect 420288 326398 420316 338014
rect 420978 337770 421006 338028
rect 421392 338014 421452 338042
rect 421576 338014 421820 338042
rect 421944 338014 422188 338042
rect 422496 338014 422648 338042
rect 422772 338014 423016 338042
rect 423140 338014 423476 338042
rect 423784 338014 423844 338042
rect 423968 338014 424212 338042
rect 424336 338014 424672 338042
rect 424796 338014 425040 338042
rect 425164 338014 425500 338042
rect 425624 338014 425868 338042
rect 426236 338014 426388 338042
rect 420978 337742 421052 337770
rect 420276 326392 420328 326398
rect 420276 326334 420328 326340
rect 420920 326392 420972 326398
rect 420920 326334 420972 326340
rect 419816 319252 419868 319258
rect 419816 319194 419868 319200
rect 419724 12096 419776 12102
rect 419724 12038 419776 12044
rect 419632 4888 419684 4894
rect 419632 4830 419684 4836
rect 420932 4826 420960 326334
rect 421024 12034 421052 337742
rect 421392 335850 421420 338014
rect 421380 335844 421432 335850
rect 421380 335786 421432 335792
rect 421576 326398 421604 338014
rect 421564 326392 421616 326398
rect 421564 326334 421616 326340
rect 421944 316034 421972 338014
rect 422496 328454 422524 338014
rect 422772 335354 422800 338014
rect 422404 328426 422524 328454
rect 422588 335326 422800 335354
rect 422300 326392 422352 326398
rect 422300 326334 422352 326340
rect 421116 316006 421972 316034
rect 421012 12028 421064 12034
rect 421012 11970 421064 11976
rect 421116 11966 421144 316006
rect 421104 11960 421156 11966
rect 421104 11902 421156 11908
rect 422312 9450 422340 326334
rect 422404 323762 422432 328426
rect 422404 323734 422524 323762
rect 422392 323604 422444 323610
rect 422392 323546 422444 323552
rect 422404 11898 422432 323546
rect 422496 13190 422524 323734
rect 422588 323610 422616 335326
rect 423140 326398 423168 338014
rect 423784 335714 423812 338014
rect 423772 335708 423824 335714
rect 423772 335650 423824 335656
rect 423128 326392 423180 326398
rect 423128 326334 423180 326340
rect 422576 323604 422628 323610
rect 422576 323546 422628 323552
rect 423680 322516 423732 322522
rect 423680 322458 423732 322464
rect 422484 13184 422536 13190
rect 422484 13126 422536 13132
rect 422392 11892 422444 11898
rect 422392 11834 422444 11840
rect 422300 9444 422352 9450
rect 422300 9386 422352 9392
rect 420184 4820 420236 4826
rect 420184 4762 420236 4768
rect 420920 4820 420972 4826
rect 420920 4762 420972 4768
rect 419540 3800 419592 3806
rect 419540 3742 419592 3748
rect 420196 480 420224 4762
rect 421380 4548 421432 4554
rect 421380 4490 421432 4496
rect 421392 480 421420 4490
rect 423692 3670 423720 322458
rect 423772 322108 423824 322114
rect 423772 322050 423824 322056
rect 423784 9382 423812 322050
rect 423968 316034 423996 338014
rect 424336 322114 424364 338014
rect 424796 322522 424824 338014
rect 425060 323468 425112 323474
rect 425060 323410 425112 323416
rect 424784 322516 424836 322522
rect 424784 322458 424836 322464
rect 424324 322108 424376 322114
rect 424324 322050 424376 322056
rect 423876 316006 423996 316034
rect 423876 11830 423904 316006
rect 423864 11824 423916 11830
rect 423864 11766 423916 11772
rect 423772 9376 423824 9382
rect 423772 9318 423824 9324
rect 425072 9314 425100 323410
rect 425164 11762 425192 338014
rect 425624 323474 425652 338014
rect 426360 335986 426388 338014
rect 426636 338014 426696 338042
rect 426820 338014 427064 338042
rect 427188 338014 427524 338042
rect 426440 336728 426492 336734
rect 426440 336670 426492 336676
rect 426348 335980 426400 335986
rect 426348 335922 426400 335928
rect 425612 323468 425664 323474
rect 425612 323410 425664 323416
rect 425152 11756 425204 11762
rect 425152 11698 425204 11704
rect 425060 9308 425112 9314
rect 425060 9250 425112 9256
rect 424968 6384 425020 6390
rect 424968 6326 425020 6332
rect 423772 4616 423824 4622
rect 423772 4558 423824 4564
rect 423680 3664 423732 3670
rect 423680 3606 423732 3612
rect 422576 3596 422628 3602
rect 422576 3538 422628 3544
rect 422588 480 422616 3538
rect 423784 480 423812 4558
rect 424980 480 425008 6326
rect 426452 3602 426480 336670
rect 426636 336462 426664 338014
rect 426624 336456 426676 336462
rect 426624 336398 426676 336404
rect 426820 316034 426848 338014
rect 427188 336734 427216 338014
rect 427878 337770 427906 338028
rect 428016 338014 428352 338042
rect 428660 338014 428720 338042
rect 428844 338014 429088 338042
rect 429304 338014 429548 338042
rect 429672 338014 429916 338042
rect 430040 338014 430376 338042
rect 427878 337742 427952 337770
rect 427176 336728 427228 336734
rect 427176 336670 427228 336676
rect 427820 330540 427872 330546
rect 427820 330482 427872 330488
rect 426544 316006 426848 316034
rect 426544 9246 426572 316006
rect 426532 9240 426584 9246
rect 426532 9182 426584 9188
rect 427268 6316 427320 6322
rect 427268 6258 427320 6264
rect 426440 3596 426492 3602
rect 426440 3538 426492 3544
rect 426164 3528 426216 3534
rect 426164 3470 426216 3476
rect 426176 480 426204 3470
rect 427280 480 427308 6258
rect 427832 5778 427860 330482
rect 427924 6390 427952 337742
rect 428016 9178 428044 338014
rect 428660 336734 428688 338014
rect 428648 336728 428700 336734
rect 428648 336670 428700 336676
rect 428844 330546 428872 338014
rect 428832 330540 428884 330546
rect 428832 330482 428884 330488
rect 429200 330540 429252 330546
rect 429200 330482 429252 330488
rect 428004 9172 428056 9178
rect 428004 9114 428056 9120
rect 427912 6384 427964 6390
rect 427912 6326 427964 6332
rect 429212 6322 429240 330482
rect 429304 9110 429332 338014
rect 429672 316034 429700 338014
rect 430040 330546 430068 338014
rect 430730 337770 430758 338028
rect 431052 338014 431112 338042
rect 431236 338014 431572 338042
rect 431696 338014 431940 338042
rect 432064 338014 432400 338042
rect 432524 338014 432768 338042
rect 432892 338014 433136 338042
rect 433536 338014 433596 338042
rect 433720 338014 433964 338042
rect 434424 338014 434668 338042
rect 434792 338014 435128 338042
rect 430730 337742 430804 337770
rect 430028 330540 430080 330546
rect 430028 330482 430080 330488
rect 430580 330540 430632 330546
rect 430580 330482 430632 330488
rect 429396 316006 429700 316034
rect 429396 13122 429424 316006
rect 429384 13116 429436 13122
rect 429384 13058 429436 13064
rect 429292 9104 429344 9110
rect 429292 9046 429344 9052
rect 429200 6316 429252 6322
rect 429200 6258 429252 6264
rect 430592 6254 430620 330482
rect 430672 330472 430724 330478
rect 430672 330414 430724 330420
rect 430684 8974 430712 330414
rect 430776 9042 430804 337742
rect 431052 335782 431080 338014
rect 431040 335776 431092 335782
rect 431040 335718 431092 335724
rect 431236 330546 431264 338014
rect 431224 330540 431276 330546
rect 431224 330482 431276 330488
rect 431696 330478 431724 338014
rect 432064 336682 432092 338014
rect 431972 336654 432092 336682
rect 431684 330472 431736 330478
rect 431684 330414 431736 330420
rect 430764 9036 430816 9042
rect 430764 8978 430816 8984
rect 430672 8968 430724 8974
rect 430672 8910 430724 8916
rect 428464 6248 428516 6254
rect 428464 6190 428516 6196
rect 430580 6248 430632 6254
rect 430580 6190 430632 6196
rect 427820 5772 427872 5778
rect 427820 5714 427872 5720
rect 428476 480 428504 6190
rect 430856 5908 430908 5914
rect 430856 5850 430908 5856
rect 429660 3460 429712 3466
rect 429660 3402 429712 3408
rect 429672 480 429700 3402
rect 430868 480 430896 5850
rect 431972 3534 432000 336654
rect 432524 335354 432552 338014
rect 432064 335326 432552 335354
rect 432064 6186 432092 335326
rect 432892 316034 432920 338014
rect 433536 336666 433564 338014
rect 433524 336660 433576 336666
rect 433524 336602 433576 336608
rect 433720 316034 433748 338014
rect 434640 336598 434668 338014
rect 434628 336592 434680 336598
rect 434628 336534 434680 336540
rect 433984 336524 434036 336530
rect 433984 336466 434036 336472
rect 432156 316006 432920 316034
rect 433352 316006 433748 316034
rect 432156 8945 432184 316006
rect 432142 8936 432198 8945
rect 432142 8871 432198 8880
rect 432052 6180 432104 6186
rect 432052 6122 432104 6128
rect 432052 5840 432104 5846
rect 432052 5782 432104 5788
rect 431960 3528 432012 3534
rect 431960 3470 432012 3476
rect 432064 480 432092 5782
rect 433248 3936 433300 3942
rect 433248 3878 433300 3884
rect 433260 480 433288 3878
rect 433352 3466 433380 316006
rect 433996 6914 434024 336466
rect 435100 336025 435128 338014
rect 435086 336016 435142 336025
rect 435086 335951 435142 335960
rect 434076 335912 434128 335918
rect 434076 335854 434128 335860
rect 433904 6886 434024 6914
rect 433904 3942 433932 6886
rect 434088 6526 434116 335854
rect 436756 16574 436784 499967
rect 577320 498704 577372 498710
rect 577320 498646 577372 498652
rect 574742 498536 574798 498545
rect 574742 498471 574798 498480
rect 451924 336728 451976 336734
rect 451924 336670 451976 336676
rect 447784 335980 447836 335986
rect 447784 335922 447836 335928
rect 440884 335844 440936 335850
rect 440884 335786 440936 335792
rect 436756 16546 436876 16574
rect 435548 8764 435600 8770
rect 435548 8706 435600 8712
rect 433984 6520 434036 6526
rect 433984 6462 434036 6468
rect 434076 6520 434128 6526
rect 434076 6462 434128 6468
rect 433892 3936 433944 3942
rect 433892 3878 433944 3884
rect 433340 3460 433392 3466
rect 433340 3402 433392 3408
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 6462
rect 435560 480 435588 8706
rect 436744 6384 436796 6390
rect 436744 6326 436796 6332
rect 436756 5778 436784 6326
rect 436744 5772 436796 5778
rect 436744 5714 436796 5720
rect 436848 5681 436876 16546
rect 439136 8832 439188 8838
rect 439136 8774 439188 8780
rect 437940 5976 437992 5982
rect 437940 5918 437992 5924
rect 436834 5672 436890 5681
rect 436834 5607 436890 5616
rect 436744 3732 436796 3738
rect 436744 3674 436796 3680
rect 436756 480 436784 3674
rect 437952 480 437980 5918
rect 439148 480 439176 8774
rect 440332 4140 440384 4146
rect 440332 4082 440384 4088
rect 440344 480 440372 4082
rect 440896 3398 440924 335786
rect 440976 335708 441028 335714
rect 440976 335650 441028 335656
rect 440988 4146 441016 335650
rect 446220 9648 446272 9654
rect 446220 9590 446272 9596
rect 442632 8900 442684 8906
rect 442632 8842 442684 8848
rect 441528 6044 441580 6050
rect 441528 5986 441580 5992
rect 440976 4140 441028 4146
rect 440976 4082 441028 4088
rect 440884 3392 440936 3398
rect 440884 3334 440936 3340
rect 441540 480 441568 5986
rect 442644 480 442672 8842
rect 445024 6112 445076 6118
rect 445024 6054 445076 6060
rect 443826 3360 443882 3369
rect 443826 3295 443882 3304
rect 443840 480 443868 3295
rect 445036 480 445064 6054
rect 446232 480 446260 9590
rect 447796 4078 447824 335922
rect 450544 335776 450596 335782
rect 450544 335718 450596 335724
rect 449808 9580 449860 9586
rect 449808 9522 449860 9528
rect 448612 6860 448664 6866
rect 448612 6802 448664 6808
rect 447416 4072 447468 4078
rect 447416 4014 447468 4020
rect 447784 4072 447836 4078
rect 447784 4014 447836 4020
rect 447428 480 447456 4014
rect 448624 480 448652 6802
rect 449820 480 449848 9522
rect 450556 3738 450584 335718
rect 451936 3942 451964 336670
rect 458824 336660 458876 336666
rect 458824 336602 458876 336608
rect 454040 12980 454092 12986
rect 454040 12922 454092 12928
rect 453304 9512 453356 9518
rect 453304 9454 453356 9460
rect 452108 6792 452160 6798
rect 452108 6734 452160 6740
rect 450912 3936 450964 3942
rect 450912 3878 450964 3884
rect 451924 3936 451976 3942
rect 451924 3878 451976 3884
rect 450544 3732 450596 3738
rect 450544 3674 450596 3680
rect 450924 480 450952 3878
rect 452120 480 452148 6734
rect 453316 480 453344 9454
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 434414 -960 434526 326
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 12922
rect 456892 10192 456944 10198
rect 456892 10134 456944 10140
rect 455696 6724 455748 6730
rect 455696 6666 455748 6672
rect 455708 480 455736 6666
rect 456904 480 456932 10134
rect 458836 3874 458864 336602
rect 472624 336592 472676 336598
rect 472624 336534 472676 336540
rect 460204 336388 460256 336394
rect 460204 336330 460256 336336
rect 459928 10260 459980 10266
rect 459928 10202 459980 10208
rect 459192 6656 459244 6662
rect 459192 6598 459244 6604
rect 458088 3868 458140 3874
rect 458088 3810 458140 3816
rect 458824 3868 458876 3874
rect 458824 3810 458876 3816
rect 458100 480 458128 3810
rect 459204 480 459232 6598
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 10202
rect 460216 3262 460244 336330
rect 460940 336320 460992 336326
rect 460940 336262 460992 336268
rect 460952 16574 460980 336262
rect 468484 336252 468536 336258
rect 468484 336194 468536 336200
rect 465724 336184 465776 336190
rect 465724 336126 465776 336132
rect 460952 16546 461624 16574
rect 460204 3256 460256 3262
rect 460204 3198 460256 3204
rect 461596 480 461624 16546
rect 465632 11552 465684 11558
rect 465632 11494 465684 11500
rect 463976 11008 464028 11014
rect 463976 10950 464028 10956
rect 462780 6588 462832 6594
rect 462780 6530 462832 6536
rect 462792 480 462820 6530
rect 463988 480 464016 10950
rect 465172 3256 465224 3262
rect 465172 3198 465224 3204
rect 465184 480 465212 3198
rect 465644 490 465672 11494
rect 465736 3126 465764 336126
rect 467472 10940 467524 10946
rect 467472 10882 467524 10888
rect 465724 3120 465776 3126
rect 465724 3062 465776 3068
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465644 462 465856 490
rect 467484 480 467512 10882
rect 468496 3194 468524 336194
rect 469862 336016 469918 336025
rect 469862 335951 469918 335960
rect 469876 16574 469904 335951
rect 469876 16546 469996 16574
rect 469864 11620 469916 11626
rect 469864 11562 469916 11568
rect 468484 3188 468536 3194
rect 468484 3130 468536 3136
rect 468668 3120 468720 3126
rect 468668 3062 468720 3068
rect 468680 480 468708 3062
rect 469876 480 469904 11562
rect 469968 3369 469996 16546
rect 470600 10872 470652 10878
rect 470600 10814 470652 10820
rect 469954 3360 470010 3369
rect 469954 3295 470010 3304
rect 465828 354 465856 462
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 10814
rect 472636 4010 472664 336534
rect 475384 336456 475436 336462
rect 475384 336398 475436 336404
rect 473452 11688 473504 11694
rect 473452 11630 473504 11636
rect 472256 4004 472308 4010
rect 472256 3946 472308 3952
rect 472624 4004 472676 4010
rect 472624 3946 472676 3952
rect 472268 480 472296 3946
rect 473464 480 473492 11630
rect 474096 10804 474148 10810
rect 474096 10746 474148 10752
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 10746
rect 475396 3262 475424 336398
rect 528560 336116 528612 336122
rect 528560 336058 528612 336064
rect 497096 13796 497148 13802
rect 497096 13738 497148 13744
rect 493048 13048 493100 13054
rect 493048 12990 493100 12996
rect 476488 12436 476540 12442
rect 476488 12378 476540 12384
rect 475752 3324 475804 3330
rect 475752 3266 475804 3272
rect 475384 3256 475436 3262
rect 475384 3198 475436 3204
rect 475764 480 475792 3266
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 12378
rect 481732 12368 481784 12374
rect 481732 12310 481784 12316
rect 478144 10736 478196 10742
rect 478144 10678 478196 10684
rect 478156 480 478184 10678
rect 480536 10600 480588 10606
rect 480536 10542 480588 10548
rect 479340 3188 479392 3194
rect 479340 3130 479392 3136
rect 479352 480 479380 3130
rect 480548 480 480576 10542
rect 481744 480 481772 12310
rect 489920 12300 489972 12306
rect 489920 12242 489972 12248
rect 482376 10668 482428 10674
rect 482376 10610 482428 10616
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 10610
rect 484032 10532 484084 10538
rect 484032 10474 484084 10480
rect 484044 480 484072 10474
rect 486424 10464 486476 10470
rect 486424 10406 486476 10412
rect 485228 7404 485280 7410
rect 485228 7346 485280 7352
rect 485240 480 485268 7346
rect 486436 480 486464 10406
rect 487160 10396 487212 10402
rect 487160 10338 487212 10344
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 10338
rect 488816 7472 488868 7478
rect 488816 7414 488868 7420
rect 488828 480 488856 7414
rect 489932 480 489960 12242
rect 490656 10328 490708 10334
rect 490656 10270 490708 10276
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 10270
rect 492312 7540 492364 7546
rect 492312 7482 492364 7488
rect 492324 480 492352 7482
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 12990
rect 494704 12232 494756 12238
rect 494704 12174 494756 12180
rect 494716 480 494744 12174
rect 495900 8288 495952 8294
rect 495900 8230 495952 8236
rect 495912 480 495940 8230
rect 497108 480 497136 13738
rect 500592 13728 500644 13734
rect 500592 13670 500644 13676
rect 499396 8220 499448 8226
rect 499396 8162 499448 8168
rect 498200 4684 498252 4690
rect 498200 4626 498252 4632
rect 498212 480 498240 4626
rect 499408 480 499436 8162
rect 500604 480 500632 13670
rect 503720 13660 503772 13666
rect 503720 13602 503772 13608
rect 502984 8152 503036 8158
rect 502984 8094 503036 8100
rect 501788 4752 501840 4758
rect 501788 4694 501840 4700
rect 501800 480 501828 4694
rect 502996 480 503024 8094
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 13602
rect 507216 13592 507268 13598
rect 507216 13534 507268 13540
rect 506480 8084 506532 8090
rect 506480 8026 506532 8032
rect 505376 5500 505428 5506
rect 505376 5442 505428 5448
rect 505388 480 505416 5442
rect 506492 480 506520 8026
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 13534
rect 511264 13524 511316 13530
rect 511264 13466 511316 13472
rect 510068 8016 510120 8022
rect 510068 7958 510120 7964
rect 508872 5432 508924 5438
rect 508872 5374 508924 5380
rect 508884 480 508912 5374
rect 510080 480 510108 7958
rect 511276 480 511304 13466
rect 514760 13456 514812 13462
rect 514760 13398 514812 13404
rect 513564 7948 513616 7954
rect 513564 7890 513616 7896
rect 512460 5364 512512 5370
rect 512460 5306 512512 5312
rect 512472 480 512500 5306
rect 513576 480 513604 7890
rect 514772 480 514800 13398
rect 521660 13388 521712 13394
rect 521660 13330 521712 13336
rect 517152 7880 517204 7886
rect 517152 7822 517204 7828
rect 515956 5296 516008 5302
rect 515956 5238 516008 5244
rect 515968 480 515996 5238
rect 517164 480 517192 7822
rect 520740 7812 520792 7818
rect 520740 7754 520792 7760
rect 518348 6520 518400 6526
rect 518348 6462 518400 6468
rect 518360 480 518388 6462
rect 519544 5228 519596 5234
rect 519544 5170 519596 5176
rect 519556 480 519584 5170
rect 520752 480 520780 7754
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521672 354 521700 13330
rect 525432 13320 525484 13326
rect 525432 13262 525484 13268
rect 524236 7744 524288 7750
rect 524236 7686 524288 7692
rect 523040 5160 523092 5166
rect 523040 5102 523092 5108
rect 523052 480 523080 5102
rect 524248 480 524276 7686
rect 525444 480 525472 13262
rect 527824 7676 527876 7682
rect 527824 7618 527876 7624
rect 526628 5092 526680 5098
rect 526628 5034 526680 5040
rect 526640 480 526668 5034
rect 527836 480 527864 7618
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 336058
rect 535460 336048 535512 336054
rect 535460 335990 535512 335996
rect 535472 16574 535500 335990
rect 574756 60722 574784 498471
rect 574836 498364 574888 498370
rect 574836 498306 574888 498312
rect 574848 100706 574876 498306
rect 577332 325514 577360 498646
rect 577412 498636 577464 498642
rect 577412 498578 577464 498584
rect 577320 325508 577372 325514
rect 577320 325450 577372 325456
rect 577424 299470 577452 498578
rect 577964 498500 578016 498506
rect 577964 498442 578016 498448
rect 577780 498432 577832 498438
rect 577594 498400 577650 498409
rect 577780 498374 577832 498380
rect 577594 498335 577650 498344
rect 577504 498228 577556 498234
rect 577504 498170 577556 498176
rect 577412 299464 577464 299470
rect 577412 299406 577464 299412
rect 577516 113014 577544 498170
rect 577504 113008 577556 113014
rect 577504 112950 577556 112956
rect 574836 100700 574888 100706
rect 574836 100642 574888 100648
rect 577608 73166 577636 498335
rect 577688 498296 577740 498302
rect 577688 498238 577740 498244
rect 577700 153202 577728 498238
rect 577792 193186 577820 498374
rect 577870 497176 577926 497185
rect 577870 497111 577926 497120
rect 577884 206990 577912 497111
rect 577976 233238 578004 498442
rect 578068 245614 578096 500142
rect 578148 498568 578200 498574
rect 578148 498510 578200 498516
rect 578160 273222 578188 498510
rect 578148 273216 578200 273222
rect 578148 273158 578200 273164
rect 578056 245608 578108 245614
rect 578056 245550 578108 245556
rect 577964 233232 578016 233238
rect 577964 233174 578016 233180
rect 577872 206984 577924 206990
rect 577872 206926 577924 206932
rect 577780 193180 577832 193186
rect 577780 193122 577832 193128
rect 577688 153196 577740 153202
rect 577688 153138 577740 153144
rect 578896 139369 578924 501026
rect 578988 179217 579016 501094
rect 579080 219065 579108 501162
rect 579172 258913 579200 502318
rect 579264 312089 579292 502386
rect 580908 498772 580960 498778
rect 580908 498714 580960 498720
rect 580172 497344 580224 497350
rect 580172 497286 580224 497292
rect 580080 497276 580132 497282
rect 580080 497218 580132 497224
rect 580092 484673 580120 497218
rect 580078 484664 580134 484673
rect 580078 484599 580134 484608
rect 580184 471481 580212 497286
rect 580724 497208 580776 497214
rect 580724 497150 580776 497156
rect 580632 497072 580684 497078
rect 580262 497040 580318 497049
rect 580632 497014 580684 497020
rect 580262 496975 580318 496984
rect 580448 497004 580500 497010
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 579250 312080 579306 312089
rect 579250 312015 579306 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 579158 258904 579214 258913
rect 579158 258839 579214 258848
rect 579620 245608 579672 245614
rect 579618 245576 579620 245585
rect 579672 245576 579674 245585
rect 579618 245511 579674 245520
rect 579804 233232 579856 233238
rect 579804 233174 579856 233180
rect 579816 232393 579844 233174
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579066 219056 579122 219065
rect 579066 218991 579122 219000
rect 579988 206984 580040 206990
rect 579988 206926 580040 206932
rect 580000 205737 580028 206926
rect 579986 205728 580042 205737
rect 579986 205663 580042 205672
rect 579620 193180 579672 193186
rect 579620 193122 579672 193128
rect 579632 192545 579660 193122
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 578974 179208 579030 179217
rect 578974 179143 579030 179152
rect 580276 165889 580304 496975
rect 580448 496946 580500 496952
rect 580356 496868 580408 496874
rect 580356 496810 580408 496816
rect 580368 351937 580396 496810
rect 580460 365129 580488 496946
rect 580540 496936 580592 496942
rect 580540 496878 580592 496884
rect 580552 378457 580580 496878
rect 580644 404977 580672 497014
rect 580736 418305 580764 497150
rect 580816 497140 580868 497146
rect 580816 497082 580868 497088
rect 580828 431633 580856 497082
rect 580920 458153 580948 498714
rect 580906 458144 580962 458153
rect 580906 458079 580962 458088
rect 580814 431624 580870 431633
rect 580814 431559 580870 431568
rect 580722 418296 580778 418305
rect 580722 418231 580778 418240
rect 580630 404968 580686 404977
rect 580630 404903 580686 404912
rect 580538 378448 580594 378457
rect 580538 378383 580594 378392
rect 580446 365120 580502 365129
rect 580446 365055 580502 365064
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580448 325508 580500 325514
rect 580448 325450 580500 325456
rect 580460 325281 580488 325450
rect 580446 325272 580502 325281
rect 580446 325207 580502 325216
rect 580262 165880 580318 165889
rect 580262 165815 580318 165824
rect 580632 153196 580684 153202
rect 580632 153138 580684 153144
rect 580644 152697 580672 153138
rect 580630 152688 580686 152697
rect 580630 152623 580686 152632
rect 578882 139360 578938 139369
rect 578882 139295 578938 139304
rect 580356 113008 580408 113014
rect 580356 112950 580408 112956
rect 580368 112849 580396 112950
rect 580354 112840 580410 112849
rect 580354 112775 580410 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 577596 73160 577648 73166
rect 577596 73102 577648 73108
rect 579712 73160 579764 73166
rect 579712 73102 579764 73108
rect 579724 73001 579752 73102
rect 579710 72992 579766 73001
rect 579710 72927 579766 72936
rect 574744 60716 574796 60722
rect 574744 60658 574796 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 535472 16546 536144 16574
rect 532056 13252 532108 13258
rect 532056 13194 532108 13200
rect 531320 7608 531372 7614
rect 531320 7550 531372 7556
rect 530124 5024 530176 5030
rect 530124 4966 530176 4972
rect 530136 480 530164 4966
rect 531332 480 531360 7550
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 354 532096 13194
rect 534448 12164 534500 12170
rect 534448 12106 534500 12112
rect 533710 4856 533766 4865
rect 533710 4791 533766 4800
rect 533724 480 533752 4791
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 12106
rect 536116 480 536144 16546
rect 546500 13184 546552 13190
rect 546500 13126 546552 13132
rect 538220 12096 538272 12102
rect 538220 12038 538272 12044
rect 537208 4956 537260 4962
rect 537208 4898 537260 4904
rect 537220 480 537248 4898
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 12038
rect 541992 12028 542044 12034
rect 541992 11970 542044 11976
rect 540796 4888 540848 4894
rect 540796 4830 540848 4836
rect 539600 3800 539652 3806
rect 539600 3742 539652 3748
rect 539612 480 539640 3742
rect 540808 480 540836 4830
rect 542004 480 542032 11970
rect 545488 11960 545540 11966
rect 545488 11902 545540 11908
rect 544384 4820 544436 4826
rect 544384 4762 544436 4768
rect 543188 3392 543240 3398
rect 543188 3334 543240 3340
rect 543200 480 543228 3334
rect 544396 480 544424 4762
rect 545500 480 545528 11902
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 13126
rect 567568 13116 567620 13122
rect 567568 13058 567620 13064
rect 547880 11892 547932 11898
rect 547880 11834 547932 11840
rect 547892 480 547920 11834
rect 551008 11824 551060 11830
rect 551008 11766 551060 11772
rect 549076 9444 549128 9450
rect 549076 9386 549128 9392
rect 549088 480 549116 9386
rect 550272 4140 550324 4146
rect 550272 4082 550324 4088
rect 550284 480 550312 4082
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 11766
rect 554780 11756 554832 11762
rect 554780 11698 554832 11704
rect 552664 9376 552716 9382
rect 552664 9318 552716 9324
rect 552676 480 552704 9318
rect 553768 3664 553820 3670
rect 553768 3606 553820 3612
rect 553780 480 553808 3606
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 11698
rect 556160 9308 556212 9314
rect 556160 9250 556212 9256
rect 556172 480 556200 9250
rect 559748 9240 559800 9246
rect 559748 9182 559800 9188
rect 557356 4072 557408 4078
rect 557356 4014 557408 4020
rect 557368 480 557396 4014
rect 558552 3324 558604 3330
rect 558552 3266 558604 3272
rect 558564 480 558592 3266
rect 559760 480 559788 9182
rect 563244 9172 563296 9178
rect 563244 9114 563296 9120
rect 562048 6452 562100 6458
rect 562048 6394 562100 6400
rect 560852 3596 560904 3602
rect 560852 3538 560904 3544
rect 560864 480 560892 3538
rect 562060 480 562088 6394
rect 563256 480 563284 9114
rect 566832 9104 566884 9110
rect 566832 9046 566884 9052
rect 565636 6384 565688 6390
rect 565636 6326 565688 6332
rect 564440 3936 564492 3942
rect 564440 3878 564492 3884
rect 564452 480 564480 3878
rect 565648 480 565676 6326
rect 566844 480 566872 9046
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 13058
rect 570328 9036 570380 9042
rect 570328 8978 570380 8984
rect 569132 6316 569184 6322
rect 569132 6258 569184 6264
rect 569144 480 569172 6258
rect 570340 480 570368 8978
rect 573916 8968 573968 8974
rect 573916 8910 573968 8916
rect 577410 8936 577466 8945
rect 572720 6248 572772 6254
rect 572720 6190 572772 6196
rect 571524 3732 571576 3738
rect 571524 3674 571576 3680
rect 571536 480 571564 3674
rect 572732 480 572760 6190
rect 573928 480 573956 8910
rect 577410 8871 577466 8880
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 575112 3528 575164 3534
rect 575112 3470 575164 3476
rect 575124 480 575152 3470
rect 576320 480 576348 6122
rect 577424 480 577452 8871
rect 582196 4004 582248 4010
rect 582196 3946 582248 3952
rect 578608 3868 578660 3874
rect 578608 3810 578660 3816
rect 578620 480 578648 3810
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3946
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 500384 3478 500440
rect 3238 475632 3294 475688
rect 3330 462576 3386 462632
rect 3054 293120 3110 293176
rect 3146 254088 3202 254144
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 4066 449520 4122 449576
rect 3974 423544 4030 423600
rect 3882 410488 3938 410544
rect 3790 397432 3846 397488
rect 3698 371320 3754 371376
rect 3606 358400 3662 358456
rect 3514 345344 3570 345400
rect 3514 306176 3570 306232
rect 3514 241032 3570 241088
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 9678 18536 9734 18592
rect 3422 6432 3478 6488
rect 5262 3304 5318 3360
rect 13542 11600 13598 11656
rect 22558 14456 22614 14512
rect 17958 12960 18014 13016
rect 140778 17176 140834 17232
rect 72606 10240 72662 10296
rect 134154 8880 134210 8936
rect 166078 7520 166134 7576
rect 233974 498752 234030 498808
rect 233882 497256 233938 497312
rect 233790 496168 233846 496224
rect 234066 497528 234122 497584
rect 235906 499976 235962 500032
rect 246670 499840 246726 499896
rect 241242 499704 241298 499760
rect 239356 498208 239412 498264
rect 244922 498480 244978 498536
rect 242806 498344 242862 498400
rect 431958 500384 432014 500440
rect 398838 500248 398894 500304
rect 403898 500112 403954 500168
rect 416226 498752 416282 498808
rect 421470 498616 421526 498672
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 436742 499976 436798 500032
rect 400494 497528 400550 497584
rect 418158 497528 418214 497584
rect 237930 497392 237986 497448
rect 251914 497392 251970 497448
rect 257158 497392 257214 497448
rect 262310 497392 262366 497448
rect 414478 497392 414534 497448
rect 419722 497392 419778 497448
rect 423862 497392 423918 497448
rect 425150 497392 425206 497448
rect 426714 497392 426770 497448
rect 428462 497392 428518 497448
rect 430210 497392 430266 497448
rect 433706 497392 433762 497448
rect 235078 496032 235134 496088
rect 200302 4800 200358 4856
rect 232226 6160 232282 6216
rect 236182 3304 236238 3360
rect 237562 18536 237618 18592
rect 240230 12960 240286 13016
rect 239034 11600 239090 11656
rect 241794 14456 241850 14512
rect 244094 3304 244150 3360
rect 259458 10240 259514 10296
rect 280250 8880 280306 8936
rect 283194 17176 283250 17232
rect 291290 7520 291346 7576
rect 296718 335960 296774 336016
rect 303710 4800 303766 4856
rect 314934 6160 314990 6216
rect 317510 3304 317566 3360
rect 336738 335960 336794 336016
rect 377862 335960 377918 336016
rect 386786 3304 386842 3360
rect 409142 335960 409198 336016
rect 416870 4800 416926 4856
rect 432142 8880 432198 8936
rect 435086 335960 435142 336016
rect 574742 498480 574798 498536
rect 436834 5616 436890 5672
rect 443826 3304 443882 3360
rect 469862 335960 469918 336016
rect 469954 3304 470010 3360
rect 577594 498344 577650 498400
rect 577870 497120 577926 497176
rect 580078 484608 580134 484664
rect 580262 496984 580318 497040
rect 580170 471416 580226 471472
rect 579250 312024 579306 312080
rect 579618 298696 579674 298752
rect 579894 272176 579950 272232
rect 579158 258848 579214 258904
rect 579618 245556 579620 245576
rect 579620 245556 579672 245576
rect 579672 245556 579674 245576
rect 579618 245520 579674 245556
rect 579802 232328 579858 232384
rect 579066 219000 579122 219056
rect 579986 205672 580042 205728
rect 579618 192480 579674 192536
rect 578974 179152 579030 179208
rect 580906 458088 580962 458144
rect 580814 431568 580870 431624
rect 580722 418240 580778 418296
rect 580630 404912 580686 404968
rect 580538 378392 580594 378448
rect 580446 365064 580502 365120
rect 580354 351872 580410 351928
rect 580446 325216 580502 325272
rect 580262 165824 580318 165880
rect 580630 152632 580686 152688
rect 578882 139304 578938 139360
rect 580354 112784 580410 112840
rect 580170 99456 580226 99512
rect 579710 72936 579766 72992
rect 580170 59608 580226 59664
rect 533710 4800 533766 4856
rect 577410 8880 577466 8936
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 3417 500442 3483 500445
rect 431953 500442 432019 500445
rect 3417 500440 432019 500442
rect 3417 500384 3422 500440
rect 3478 500384 431958 500440
rect 432014 500384 432019 500440
rect 3417 500382 432019 500384
rect 3417 500379 3483 500382
rect 431953 500379 432019 500382
rect 236678 500244 236684 500308
rect 236748 500306 236754 500308
rect 398833 500306 398899 500309
rect 236748 500304 398899 500306
rect 236748 500248 398838 500304
rect 398894 500248 398899 500304
rect 236748 500246 398899 500248
rect 236748 500244 236754 500246
rect 398833 500243 398899 500246
rect 236494 500108 236500 500172
rect 236564 500170 236570 500172
rect 403893 500170 403959 500173
rect 236564 500168 403959 500170
rect 236564 500112 403898 500168
rect 403954 500112 403959 500168
rect 236564 500110 403959 500112
rect 236564 500108 236570 500110
rect 403893 500107 403959 500110
rect 235901 500034 235967 500037
rect 436737 500034 436803 500037
rect 235901 500032 436803 500034
rect 235901 499976 235906 500032
rect 235962 499976 436742 500032
rect 436798 499976 436803 500032
rect 235901 499974 436803 499976
rect 235901 499971 235967 499974
rect 436737 499971 436803 499974
rect 246665 499898 246731 499901
rect 580390 499898 580396 499900
rect 246665 499896 580396 499898
rect 246665 499840 246670 499896
rect 246726 499840 580396 499896
rect 246665 499838 580396 499840
rect 246665 499835 246731 499838
rect 580390 499836 580396 499838
rect 580460 499836 580466 499900
rect 241237 499762 241303 499765
rect 580206 499762 580212 499764
rect 241237 499760 580212 499762
rect 241237 499704 241242 499760
rect 241298 499704 580212 499760
rect 241237 499702 580212 499704
rect 241237 499699 241303 499702
rect 580206 499700 580212 499702
rect 580276 499700 580282 499764
rect 233969 498810 234035 498813
rect 416221 498810 416287 498813
rect 233969 498808 416287 498810
rect 233969 498752 233974 498808
rect 234030 498752 416226 498808
rect 416282 498752 416287 498808
rect 233969 498750 416287 498752
rect 233969 498747 234035 498750
rect 416221 498747 416287 498750
rect 233734 498612 233740 498676
rect 233804 498674 233810 498676
rect 421465 498674 421531 498677
rect 233804 498672 421531 498674
rect 233804 498616 421470 498672
rect 421526 498616 421531 498672
rect 233804 498614 421531 498616
rect 233804 498612 233810 498614
rect 421465 498611 421531 498614
rect 244917 498538 244983 498541
rect 574737 498538 574803 498541
rect 244917 498536 574803 498538
rect 244917 498480 244922 498536
rect 244978 498480 574742 498536
rect 574798 498480 574803 498536
rect 244917 498478 574803 498480
rect 244917 498475 244983 498478
rect 574737 498475 574803 498478
rect 242801 498402 242867 498405
rect 577589 498402 577655 498405
rect 242801 498400 577655 498402
rect 242801 498344 242806 498400
rect 242862 498344 577594 498400
rect 577650 498344 577655 498400
rect 242801 498342 577655 498344
rect 242801 498339 242867 498342
rect 577589 498339 577655 498342
rect 239351 498266 239417 498269
rect 577446 498266 577452 498268
rect 239351 498264 577452 498266
rect 239351 498208 239356 498264
rect 239412 498208 577452 498264
rect 239351 498206 577452 498208
rect 239351 498203 239417 498206
rect 577446 498204 577452 498206
rect 577516 498204 577522 498268
rect 583520 497844 584960 498084
rect 234061 497586 234127 497589
rect 400489 497588 400555 497589
rect 418153 497588 418219 497589
rect 400438 497586 400444 497588
rect 234061 497584 267750 497586
rect 234061 497528 234066 497584
rect 234122 497528 267750 497584
rect 234061 497526 267750 497528
rect 400398 497526 400444 497586
rect 400508 497584 400555 497588
rect 418102 497586 418108 497588
rect 400550 497528 400555 497584
rect 234061 497523 234127 497526
rect 237925 497450 237991 497453
rect 238518 497450 238524 497452
rect 237925 497448 238524 497450
rect 237925 497392 237930 497448
rect 237986 497392 238524 497448
rect 237925 497390 238524 497392
rect 237925 497387 237991 497390
rect 238518 497388 238524 497390
rect 238588 497388 238594 497452
rect 251909 497450 251975 497453
rect 254894 497450 254900 497452
rect 251909 497448 254900 497450
rect 251909 497392 251914 497448
rect 251970 497392 254900 497448
rect 251909 497390 254900 497392
rect 251909 497387 251975 497390
rect 254894 497388 254900 497390
rect 254964 497388 254970 497452
rect 257153 497450 257219 497453
rect 262070 497450 262076 497452
rect 257153 497448 262076 497450
rect 257153 497392 257158 497448
rect 257214 497392 262076 497448
rect 257153 497390 262076 497392
rect 257153 497387 257219 497390
rect 262070 497388 262076 497390
rect 262140 497388 262146 497452
rect 262305 497450 262371 497453
rect 262305 497448 264898 497450
rect 262305 497392 262310 497448
rect 262366 497392 264898 497448
rect 262305 497390 264898 497392
rect 262305 497387 262371 497390
rect 233877 497314 233943 497317
rect 264646 497314 264652 497316
rect 233877 497312 264652 497314
rect 233877 497256 233882 497312
rect 233938 497256 264652 497312
rect 233877 497254 264652 497256
rect 233877 497251 233943 497254
rect 264646 497252 264652 497254
rect 264716 497252 264722 497316
rect 264838 497178 264898 497390
rect 265014 497388 265020 497452
rect 265084 497450 265090 497452
rect 267690 497450 267750 497526
rect 400438 497524 400444 497526
rect 400508 497524 400555 497528
rect 418062 497526 418108 497586
rect 418172 497584 418219 497588
rect 418214 497528 418219 497584
rect 418102 497524 418108 497526
rect 418172 497524 418219 497528
rect 400489 497523 400555 497524
rect 418153 497523 418219 497524
rect 414473 497450 414539 497453
rect 419717 497450 419783 497453
rect 265084 497390 265266 497450
rect 267690 497448 414539 497450
rect 267690 497392 414478 497448
rect 414534 497392 414539 497448
rect 267690 497390 414539 497392
rect 265084 497388 265090 497390
rect 265206 497314 265266 497390
rect 414473 497387 414539 497390
rect 416270 497448 419783 497450
rect 416270 497392 419722 497448
rect 419778 497392 419783 497448
rect 416270 497390 419783 497392
rect 416270 497314 416330 497390
rect 419717 497387 419783 497390
rect 423857 497450 423923 497453
rect 425145 497452 425211 497453
rect 423990 497450 423996 497452
rect 423857 497448 423996 497450
rect 423857 497392 423862 497448
rect 423918 497392 423996 497448
rect 423857 497390 423996 497392
rect 423857 497387 423923 497390
rect 423990 497388 423996 497390
rect 424060 497388 424066 497452
rect 425094 497450 425100 497452
rect 425054 497390 425100 497450
rect 425164 497448 425211 497452
rect 425206 497392 425211 497448
rect 425094 497388 425100 497390
rect 425164 497388 425211 497392
rect 426382 497388 426388 497452
rect 426452 497450 426458 497452
rect 426709 497450 426775 497453
rect 426452 497448 426775 497450
rect 426452 497392 426714 497448
rect 426770 497392 426775 497448
rect 426452 497390 426775 497392
rect 426452 497388 426458 497390
rect 425145 497387 425211 497388
rect 426709 497387 426775 497390
rect 427854 497388 427860 497452
rect 427924 497450 427930 497452
rect 428457 497450 428523 497453
rect 427924 497448 428523 497450
rect 427924 497392 428462 497448
rect 428518 497392 428523 497448
rect 427924 497390 428523 497392
rect 427924 497388 427930 497390
rect 428457 497387 428523 497390
rect 429142 497388 429148 497452
rect 429212 497450 429218 497452
rect 430205 497450 430271 497453
rect 429212 497448 430271 497450
rect 429212 497392 430210 497448
rect 430266 497392 430271 497448
rect 429212 497390 430271 497392
rect 429212 497388 429218 497390
rect 430205 497387 430271 497390
rect 433374 497388 433380 497452
rect 433444 497450 433450 497452
rect 433701 497450 433767 497453
rect 433444 497448 433767 497450
rect 433444 497392 433706 497448
rect 433762 497392 433767 497448
rect 433444 497390 433767 497392
rect 433444 497388 433450 497390
rect 433701 497387 433767 497390
rect 265206 497254 416330 497314
rect 577865 497178 577931 497181
rect 264838 497176 577931 497178
rect 264838 497120 577870 497176
rect 577926 497120 577931 497176
rect 264838 497118 577931 497120
rect 577865 497115 577931 497118
rect 262070 496980 262076 497044
rect 262140 497042 262146 497044
rect 580257 497042 580323 497045
rect 262140 497040 580323 497042
rect 262140 496984 580262 497040
rect 580318 496984 580323 497040
rect 262140 496982 580323 496984
rect 262140 496980 262146 496982
rect 580257 496979 580323 496982
rect 254894 496844 254900 496908
rect 254964 496906 254970 496908
rect 580574 496906 580580 496908
rect 254964 496846 580580 496906
rect 254964 496844 254970 496846
rect 580574 496844 580580 496846
rect 580644 496844 580650 496908
rect 233785 496226 233851 496229
rect 400438 496226 400444 496228
rect 233785 496224 400444 496226
rect 233785 496168 233790 496224
rect 233846 496168 400444 496224
rect 233785 496166 400444 496168
rect 233785 496163 233851 496166
rect 400438 496164 400444 496166
rect 400508 496164 400514 496228
rect 235073 496090 235139 496093
rect 418102 496090 418108 496092
rect 235073 496088 418108 496090
rect 235073 496032 235078 496088
rect 235134 496032 418108 496088
rect 235073 496030 418108 496032
rect 235073 496027 235139 496030
rect 418102 496028 418108 496030
rect 418172 496028 418178 496092
rect -960 488596 480 488836
rect 580073 484666 580139 484669
rect 583520 484666 584960 484756
rect 580073 484664 584960 484666
rect 580073 484608 580078 484664
rect 580134 484608 584960 484664
rect 580073 484606 584960 484608
rect 580073 484603 580139 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3233 475690 3299 475693
rect -960 475688 3299 475690
rect -960 475632 3238 475688
rect 3294 475632 3299 475688
rect -960 475630 3299 475632
rect -960 475540 480 475630
rect 3233 475627 3299 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580901 458146 580967 458149
rect 583520 458146 584960 458236
rect 580901 458144 584960 458146
rect 580901 458088 580906 458144
rect 580962 458088 584960 458144
rect 580901 458086 584960 458088
rect 580901 458083 580967 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 4061 449578 4127 449581
rect -960 449576 4127 449578
rect -960 449520 4066 449576
rect 4122 449520 4127 449576
rect -960 449518 4127 449520
rect -960 449428 480 449518
rect 4061 449515 4127 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580809 431626 580875 431629
rect 583520 431626 584960 431716
rect 580809 431624 584960 431626
rect 580809 431568 580814 431624
rect 580870 431568 584960 431624
rect 580809 431566 584960 431568
rect 580809 431563 580875 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3969 423602 4035 423605
rect -960 423600 4035 423602
rect -960 423544 3974 423600
rect 4030 423544 4035 423600
rect -960 423542 4035 423544
rect -960 423452 480 423542
rect 3969 423539 4035 423542
rect 580717 418298 580783 418301
rect 583520 418298 584960 418388
rect 580717 418296 584960 418298
rect 580717 418240 580722 418296
rect 580778 418240 584960 418296
rect 580717 418238 584960 418240
rect 580717 418235 580783 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3877 410546 3943 410549
rect -960 410544 3943 410546
rect -960 410488 3882 410544
rect 3938 410488 3943 410544
rect -960 410486 3943 410488
rect -960 410396 480 410486
rect 3877 410483 3943 410486
rect 580625 404970 580691 404973
rect 583520 404970 584960 405060
rect 580625 404968 584960 404970
rect 580625 404912 580630 404968
rect 580686 404912 584960 404968
rect 580625 404910 584960 404912
rect 580625 404907 580691 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3785 397490 3851 397493
rect -960 397488 3851 397490
rect -960 397432 3790 397488
rect 3846 397432 3851 397488
rect -960 397430 3851 397432
rect -960 397340 480 397430
rect 3785 397427 3851 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580533 378450 580599 378453
rect 583520 378450 584960 378540
rect 580533 378448 584960 378450
rect 580533 378392 580538 378448
rect 580594 378392 584960 378448
rect 580533 378390 584960 378392
rect 580533 378387 580599 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3693 371378 3759 371381
rect -960 371376 3759 371378
rect -960 371320 3698 371376
rect 3754 371320 3759 371376
rect -960 371318 3759 371320
rect -960 371228 480 371318
rect 3693 371315 3759 371318
rect 580441 365122 580507 365125
rect 583520 365122 584960 365212
rect 580441 365120 584960 365122
rect 580441 365064 580446 365120
rect 580502 365064 584960 365120
rect 580441 365062 584960 365064
rect 580441 365059 580507 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 583520 338452 584960 338692
rect 296713 336018 296779 336021
rect 336733 336018 336799 336021
rect 296713 336016 336799 336018
rect 296713 335960 296718 336016
rect 296774 335960 336738 336016
rect 336794 335960 336799 336016
rect 296713 335958 336799 335960
rect 296713 335955 296779 335958
rect 336733 335955 336799 335958
rect 377857 336018 377923 336021
rect 409137 336018 409203 336021
rect 377857 336016 409203 336018
rect 377857 335960 377862 336016
rect 377918 335960 409142 336016
rect 409198 335960 409203 336016
rect 377857 335958 409203 335960
rect 377857 335955 377923 335958
rect 409137 335955 409203 335958
rect 435081 336018 435147 336021
rect 469857 336018 469923 336021
rect 435081 336016 469923 336018
rect 435081 335960 435086 336016
rect 435142 335960 469862 336016
rect 469918 335960 469923 336016
rect 435081 335958 469923 335960
rect 435081 335955 435147 335958
rect 469857 335955 469923 335958
rect -960 332196 480 332436
rect 580441 325274 580507 325277
rect 583520 325274 584960 325364
rect 580441 325272 584960 325274
rect 580441 325216 580446 325272
rect 580502 325216 584960 325272
rect 580441 325214 584960 325216
rect 580441 325211 580507 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect -960 319230 6930 319290
rect -960 319140 480 319230
rect 6870 318882 6930 319230
rect 236678 318882 236684 318884
rect 6870 318822 236684 318882
rect 236678 318820 236684 318822
rect 236748 318820 236754 318884
rect 579245 312082 579311 312085
rect 583520 312082 584960 312172
rect 579245 312080 584960 312082
rect 579245 312024 579250 312080
rect 579306 312024 584960 312080
rect 579245 312022 584960 312024
rect 579245 312019 579311 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect -960 267142 674 267202
rect -960 267066 480 267142
rect 614 267066 674 267142
rect -960 267052 674 267066
rect 246 267006 674 267052
rect 246 266522 306 267006
rect 246 266462 6930 266522
rect 6870 266386 6930 266462
rect 236494 266386 236500 266388
rect 6870 266326 236500 266386
rect 236494 266324 236500 266326
rect 236564 266324 236570 266388
rect 579153 258906 579219 258909
rect 583520 258906 584960 258996
rect 579153 258904 584960 258906
rect 579153 258848 579158 258904
rect 579214 258848 584960 258904
rect 579153 258846 584960 258848
rect 579153 258843 579219 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 579613 245578 579679 245581
rect 583520 245578 584960 245668
rect 579613 245576 584960 245578
rect 579613 245520 579618 245576
rect 579674 245520 584960 245576
rect 579613 245518 584960 245520
rect 579613 245515 579679 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579061 219058 579127 219061
rect 583520 219058 584960 219148
rect 579061 219056 584960 219058
rect 579061 219000 579066 219056
rect 579122 219000 584960 219056
rect 579061 218998 584960 219000
rect 579061 218995 579127 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579981 205730 580047 205733
rect 583520 205730 584960 205820
rect 579981 205728 584960 205730
rect 579981 205672 579986 205728
rect 580042 205672 584960 205728
rect 579981 205670 584960 205672
rect 579981 205667 580047 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 578969 179210 579035 179213
rect 583520 179210 584960 179300
rect 578969 179208 584960 179210
rect 578969 179152 578974 179208
rect 579030 179152 584960 179208
rect 578969 179150 584960 179152
rect 578969 179147 579035 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580257 165882 580323 165885
rect 583520 165882 584960 165972
rect 580257 165880 584960 165882
rect 580257 165824 580262 165880
rect 580318 165824 584960 165880
rect 580257 165822 584960 165824
rect 580257 165819 580323 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580625 152690 580691 152693
rect 583520 152690 584960 152780
rect 580625 152688 584960 152690
rect 580625 152632 580630 152688
rect 580686 152632 584960 152688
rect 580625 152630 584960 152632
rect 580625 152627 580691 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 578877 139362 578943 139365
rect 583520 139362 584960 139452
rect 578877 139360 584960 139362
rect 578877 139304 578882 139360
rect 578938 139304 584960 139360
rect 578877 139302 584960 139304
rect 578877 139299 578943 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580574 125972 580580 126036
rect 580644 126034 580650 126036
rect 583520 126034 584960 126124
rect 580644 125974 584960 126034
rect 580644 125972 580650 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580349 112842 580415 112845
rect 583520 112842 584960 112932
rect 580349 112840 584960 112842
rect 580349 112784 580354 112840
rect 580410 112784 584960 112840
rect 580349 112782 584960 112784
rect 580349 112779 580415 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect -960 97550 674 97610
rect -960 97474 480 97550
rect 614 97474 674 97550
rect -960 97460 674 97474
rect 246 97414 674 97460
rect 246 96930 306 97414
rect 246 96870 6930 96930
rect 6870 96658 6930 96870
rect 423990 96658 423996 96660
rect 6870 96598 423996 96658
rect 423990 96596 423996 96598
rect 424060 96596 424066 96660
rect 580390 86124 580396 86188
rect 580460 86186 580466 86188
rect 583520 86186 584960 86276
rect 580460 86126 584960 86186
rect 580460 86124 580466 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect -960 84630 6930 84690
rect -960 84540 480 84630
rect 6870 84282 6930 84630
rect 233734 84282 233740 84284
rect 6870 84222 233740 84282
rect 233734 84220 233740 84222
rect 233804 84220 233810 84284
rect 579705 72994 579771 72997
rect 583520 72994 584960 73084
rect 579705 72992 584960 72994
rect 579705 72936 579710 72992
rect 579766 72936 584960 72992
rect 579705 72934 584960 72936
rect 579705 72931 579771 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect -960 71574 674 71634
rect -960 71498 480 71574
rect 614 71498 674 71574
rect -960 71484 674 71498
rect 246 71438 674 71484
rect 246 70954 306 71438
rect 246 70894 6930 70954
rect 6870 70410 6930 70894
rect 425094 70410 425100 70412
rect 6870 70350 425100 70410
rect 425094 70348 425100 70350
rect 425164 70348 425170 70412
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect -960 58518 674 58578
rect -960 58442 480 58518
rect 614 58442 674 58518
rect -960 58428 674 58442
rect 246 58382 674 58428
rect 246 58034 306 58382
rect 427854 58034 427860 58036
rect 246 57974 427860 58034
rect 427854 57972 427860 57974
rect 427924 57972 427930 58036
rect 580206 46276 580212 46340
rect 580276 46338 580282 46340
rect 583520 46338 584960 46428
rect 580276 46278 584960 46338
rect 580276 46276 580282 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 426382 44298 426388 44300
rect 6870 44238 426388 44298
rect 426382 44236 426388 44238
rect 426452 44236 426458 44300
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect -960 32406 674 32466
rect -960 32330 480 32406
rect 614 32330 674 32406
rect -960 32316 674 32330
rect 246 32270 674 32316
rect 246 31786 306 32270
rect 238518 31860 238524 31924
rect 238588 31922 238594 31924
rect 583526 31922 583586 32950
rect 238588 31862 583586 31922
rect 238588 31860 238594 31862
rect 429142 31786 429148 31788
rect 246 31726 429148 31786
rect 429142 31724 429148 31726
rect 429212 31724 429218 31788
rect 577446 19756 577452 19820
rect 577516 19818 577522 19820
rect 583520 19818 584960 19908
rect 577516 19758 584960 19818
rect 577516 19756 577522 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 433374 19410 433380 19412
rect -960 19350 433380 19410
rect -960 19260 480 19350
rect 433374 19348 433380 19350
rect 433444 19348 433450 19412
rect 9673 18594 9739 18597
rect 237557 18594 237623 18597
rect 9673 18592 237623 18594
rect 9673 18536 9678 18592
rect 9734 18536 237562 18592
rect 237618 18536 237623 18592
rect 9673 18534 237623 18536
rect 9673 18531 9739 18534
rect 237557 18531 237623 18534
rect 140773 17234 140839 17237
rect 283189 17234 283255 17237
rect 140773 17232 283255 17234
rect 140773 17176 140778 17232
rect 140834 17176 283194 17232
rect 283250 17176 283255 17232
rect 140773 17174 283255 17176
rect 140773 17171 140839 17174
rect 283189 17171 283255 17174
rect 22553 14514 22619 14517
rect 241789 14514 241855 14517
rect 22553 14512 241855 14514
rect 22553 14456 22558 14512
rect 22614 14456 241794 14512
rect 241850 14456 241855 14512
rect 22553 14454 241855 14456
rect 22553 14451 22619 14454
rect 241789 14451 241855 14454
rect 17953 13018 18019 13021
rect 240225 13018 240291 13021
rect 17953 13016 240291 13018
rect 17953 12960 17958 13016
rect 18014 12960 240230 13016
rect 240286 12960 240291 13016
rect 17953 12958 240291 12960
rect 17953 12955 18019 12958
rect 240225 12955 240291 12958
rect 13537 11658 13603 11661
rect 239029 11658 239095 11661
rect 13537 11656 239095 11658
rect 13537 11600 13542 11656
rect 13598 11600 239034 11656
rect 239090 11600 239095 11656
rect 13537 11598 239095 11600
rect 13537 11595 13603 11598
rect 239029 11595 239095 11598
rect 72601 10298 72667 10301
rect 259453 10298 259519 10301
rect 72601 10296 259519 10298
rect 72601 10240 72606 10296
rect 72662 10240 259458 10296
rect 259514 10240 259519 10296
rect 72601 10238 259519 10240
rect 72601 10235 72667 10238
rect 259453 10235 259519 10238
rect 134149 8938 134215 8941
rect 280245 8938 280311 8941
rect 134149 8936 280311 8938
rect 134149 8880 134154 8936
rect 134210 8880 280250 8936
rect 280306 8880 280311 8936
rect 134149 8878 280311 8880
rect 134149 8875 134215 8878
rect 280245 8875 280311 8878
rect 432137 8938 432203 8941
rect 577405 8938 577471 8941
rect 432137 8936 577471 8938
rect 432137 8880 432142 8936
rect 432198 8880 577410 8936
rect 577466 8880 577471 8936
rect 432137 8878 577471 8880
rect 432137 8875 432203 8878
rect 577405 8875 577471 8878
rect 166073 7578 166139 7581
rect 291285 7578 291351 7581
rect 166073 7576 291351 7578
rect 166073 7520 166078 7576
rect 166134 7520 291290 7576
rect 291346 7520 291351 7576
rect 166073 7518 291351 7520
rect 166073 7515 166139 7518
rect 291285 7515 291351 7518
rect 583520 6626 584960 6716
rect -960 6490 480 6580
rect 583342 6566 584960 6626
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect 583342 6490 583402 6566
rect 583520 6490 584960 6566
rect 583342 6476 584960 6490
rect 583342 6430 583586 6476
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 232221 6218 232287 6221
rect 314929 6218 314995 6221
rect 232221 6216 314995 6218
rect 232221 6160 232226 6216
rect 232282 6160 314934 6216
rect 314990 6160 314995 6216
rect 232221 6158 314995 6160
rect 232221 6155 232287 6158
rect 314929 6155 314995 6158
rect 436829 5674 436895 5677
rect 583526 5674 583586 6430
rect 436829 5672 583586 5674
rect 436829 5616 436834 5672
rect 436890 5616 583586 5672
rect 436829 5614 583586 5616
rect 436829 5611 436895 5614
rect 200297 4858 200363 4861
rect 303705 4858 303771 4861
rect 200297 4856 303771 4858
rect 200297 4800 200302 4856
rect 200358 4800 303710 4856
rect 303766 4800 303771 4856
rect 200297 4798 303771 4800
rect 200297 4795 200363 4798
rect 303705 4795 303771 4798
rect 416865 4858 416931 4861
rect 533705 4858 533771 4861
rect 416865 4856 533771 4858
rect 416865 4800 416870 4856
rect 416926 4800 533710 4856
rect 533766 4800 533771 4856
rect 416865 4798 533771 4800
rect 416865 4795 416931 4798
rect 533705 4795 533771 4798
rect 5257 3362 5323 3365
rect 236177 3362 236243 3365
rect 5257 3360 236243 3362
rect 5257 3304 5262 3360
rect 5318 3304 236182 3360
rect 236238 3304 236243 3360
rect 5257 3302 236243 3304
rect 5257 3299 5323 3302
rect 236177 3299 236243 3302
rect 244089 3362 244155 3365
rect 317505 3362 317571 3365
rect 244089 3360 317571 3362
rect 244089 3304 244094 3360
rect 244150 3304 317510 3360
rect 317566 3304 317571 3360
rect 244089 3302 317571 3304
rect 244089 3299 244155 3302
rect 317505 3299 317571 3302
rect 386781 3362 386847 3365
rect 443821 3362 443887 3365
rect 386781 3360 443887 3362
rect 386781 3304 386786 3360
rect 386842 3304 443826 3360
rect 443882 3304 443887 3360
rect 386781 3302 443887 3304
rect 386781 3299 386847 3302
rect 443821 3299 443887 3302
rect 469949 3362 470015 3365
rect 583385 3362 583451 3365
rect 469949 3360 583451 3362
rect 469949 3304 469954 3360
rect 470010 3304 583390 3360
rect 583446 3304 583451 3360
rect 469949 3302 583451 3304
rect 469949 3299 470015 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 236684 500244 236748 500308
rect 236500 500108 236564 500172
rect 580396 499836 580460 499900
rect 580212 499700 580276 499764
rect 233740 498612 233804 498676
rect 577452 498204 577516 498268
rect 400444 497584 400508 497588
rect 400444 497528 400494 497584
rect 400494 497528 400508 497584
rect 238524 497388 238588 497452
rect 254900 497388 254964 497452
rect 262076 497388 262140 497452
rect 264652 497252 264716 497316
rect 265020 497388 265084 497452
rect 400444 497524 400508 497528
rect 418108 497584 418172 497588
rect 418108 497528 418158 497584
rect 418158 497528 418172 497584
rect 418108 497524 418172 497528
rect 423996 497388 424060 497452
rect 425100 497448 425164 497452
rect 425100 497392 425150 497448
rect 425150 497392 425164 497448
rect 425100 497388 425164 497392
rect 426388 497388 426452 497452
rect 427860 497388 427924 497452
rect 429148 497388 429212 497452
rect 433380 497388 433444 497452
rect 262076 496980 262140 497044
rect 254900 496844 254964 496908
rect 580580 496844 580644 496908
rect 400444 496164 400508 496228
rect 418108 496028 418172 496092
rect 236684 318820 236748 318884
rect 236500 266324 236564 266388
rect 580580 125972 580644 126036
rect 423996 96596 424060 96660
rect 580396 86124 580460 86188
rect 233740 84220 233804 84284
rect 425100 70348 425164 70412
rect 427860 57972 427924 58036
rect 580212 46276 580276 46340
rect 426388 44236 426452 44300
rect 238524 31860 238588 31924
rect 429148 31724 429212 31788
rect 577452 19756 577516 19820
rect 433380 19348 433444 19412
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 680614 -8106 711002
rect -8726 680058 -8694 680614
rect -8138 680058 -8106 680614
rect -8726 644614 -8106 680058
rect -8726 644058 -8694 644614
rect -8138 644058 -8106 644614
rect -8726 608614 -8106 644058
rect -8726 608058 -8694 608614
rect -8138 608058 -8106 608614
rect -8726 572614 -8106 608058
rect -8726 572058 -8694 572614
rect -8138 572058 -8106 572614
rect -8726 536614 -8106 572058
rect -8726 536058 -8694 536614
rect -8138 536058 -8106 536614
rect -8726 500614 -8106 536058
rect -8726 500058 -8694 500614
rect -8138 500058 -8106 500614
rect -8726 464614 -8106 500058
rect -8726 464058 -8694 464614
rect -8138 464058 -8106 464614
rect -8726 428614 -8106 464058
rect -8726 428058 -8694 428614
rect -8138 428058 -8106 428614
rect -8726 392614 -8106 428058
rect -8726 392058 -8694 392614
rect -8138 392058 -8106 392614
rect -8726 356614 -8106 392058
rect -8726 356058 -8694 356614
rect -8138 356058 -8106 356614
rect -8726 320614 -8106 356058
rect -8726 320058 -8694 320614
rect -8138 320058 -8106 320614
rect -8726 284614 -8106 320058
rect -8726 284058 -8694 284614
rect -8138 284058 -8106 284614
rect -8726 248614 -8106 284058
rect -8726 248058 -8694 248614
rect -8138 248058 -8106 248614
rect -8726 212614 -8106 248058
rect -8726 212058 -8694 212614
rect -8138 212058 -8106 212614
rect -8726 176614 -8106 212058
rect -8726 176058 -8694 176614
rect -8138 176058 -8106 176614
rect -8726 140614 -8106 176058
rect -8726 140058 -8694 140614
rect -8138 140058 -8106 140614
rect -8726 104614 -8106 140058
rect -8726 104058 -8694 104614
rect -8138 104058 -8106 104614
rect -8726 68614 -8106 104058
rect -8726 68058 -8694 68614
rect -8138 68058 -8106 68614
rect -8726 32614 -8106 68058
rect -8726 32058 -8694 32614
rect -8138 32058 -8106 32614
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710042 12986 710598
rect 13542 710042 13574 710598
rect -7766 698058 -7734 698614
rect -7178 698058 -7146 698614
rect -7766 662614 -7146 698058
rect -7766 662058 -7734 662614
rect -7178 662058 -7146 662614
rect -7766 626614 -7146 662058
rect -7766 626058 -7734 626614
rect -7178 626058 -7146 626614
rect -7766 590614 -7146 626058
rect -7766 590058 -7734 590614
rect -7178 590058 -7146 590614
rect -7766 554614 -7146 590058
rect -7766 554058 -7734 554614
rect -7178 554058 -7146 554614
rect -7766 518614 -7146 554058
rect -7766 518058 -7734 518614
rect -7178 518058 -7146 518614
rect -7766 482614 -7146 518058
rect -7766 482058 -7734 482614
rect -7178 482058 -7146 482614
rect -7766 446614 -7146 482058
rect -7766 446058 -7734 446614
rect -7178 446058 -7146 446614
rect -7766 410614 -7146 446058
rect -7766 410058 -7734 410614
rect -7178 410058 -7146 410614
rect -7766 374614 -7146 410058
rect -7766 374058 -7734 374614
rect -7178 374058 -7146 374614
rect -7766 338614 -7146 374058
rect -7766 338058 -7734 338614
rect -7178 338058 -7146 338614
rect -7766 302614 -7146 338058
rect -7766 302058 -7734 302614
rect -7178 302058 -7146 302614
rect -7766 266614 -7146 302058
rect -7766 266058 -7734 266614
rect -7178 266058 -7146 266614
rect -7766 230614 -7146 266058
rect -7766 230058 -7734 230614
rect -7178 230058 -7146 230614
rect -7766 194614 -7146 230058
rect -7766 194058 -7734 194614
rect -7178 194058 -7146 194614
rect -7766 158614 -7146 194058
rect -7766 158058 -7734 158614
rect -7178 158058 -7146 158614
rect -7766 122614 -7146 158058
rect -7766 122058 -7734 122614
rect -7178 122058 -7146 122614
rect -7766 86614 -7146 122058
rect -7766 86058 -7734 86614
rect -7178 86058 -7146 86614
rect -7766 50614 -7146 86058
rect -7766 50058 -7734 50614
rect -7178 50058 -7146 50614
rect -7766 14614 -7146 50058
rect -7766 14058 -7734 14614
rect -7178 14058 -7146 14614
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 676894 -6186 709082
rect -6806 676338 -6774 676894
rect -6218 676338 -6186 676894
rect -6806 640894 -6186 676338
rect -6806 640338 -6774 640894
rect -6218 640338 -6186 640894
rect -6806 604894 -6186 640338
rect -6806 604338 -6774 604894
rect -6218 604338 -6186 604894
rect -6806 568894 -6186 604338
rect -6806 568338 -6774 568894
rect -6218 568338 -6186 568894
rect -6806 532894 -6186 568338
rect -6806 532338 -6774 532894
rect -6218 532338 -6186 532894
rect -6806 496894 -6186 532338
rect -6806 496338 -6774 496894
rect -6218 496338 -6186 496894
rect -6806 460894 -6186 496338
rect -6806 460338 -6774 460894
rect -6218 460338 -6186 460894
rect -6806 424894 -6186 460338
rect -6806 424338 -6774 424894
rect -6218 424338 -6186 424894
rect -6806 388894 -6186 424338
rect -6806 388338 -6774 388894
rect -6218 388338 -6186 388894
rect -6806 352894 -6186 388338
rect -6806 352338 -6774 352894
rect -6218 352338 -6186 352894
rect -6806 316894 -6186 352338
rect -6806 316338 -6774 316894
rect -6218 316338 -6186 316894
rect -6806 280894 -6186 316338
rect -6806 280338 -6774 280894
rect -6218 280338 -6186 280894
rect -6806 244894 -6186 280338
rect -6806 244338 -6774 244894
rect -6218 244338 -6186 244894
rect -6806 208894 -6186 244338
rect -6806 208338 -6774 208894
rect -6218 208338 -6186 208894
rect -6806 172894 -6186 208338
rect -6806 172338 -6774 172894
rect -6218 172338 -6186 172894
rect -6806 136894 -6186 172338
rect -6806 136338 -6774 136894
rect -6218 136338 -6186 136894
rect -6806 100894 -6186 136338
rect -6806 100338 -6774 100894
rect -6218 100338 -6186 100894
rect -6806 64894 -6186 100338
rect -6806 64338 -6774 64894
rect -6218 64338 -6186 64894
rect -6806 28894 -6186 64338
rect -6806 28338 -6774 28894
rect -6218 28338 -6186 28894
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708122 9266 708678
rect 9822 708122 9854 708678
rect -5846 694338 -5814 694894
rect -5258 694338 -5226 694894
rect -5846 658894 -5226 694338
rect -5846 658338 -5814 658894
rect -5258 658338 -5226 658894
rect -5846 622894 -5226 658338
rect -5846 622338 -5814 622894
rect -5258 622338 -5226 622894
rect -5846 586894 -5226 622338
rect -5846 586338 -5814 586894
rect -5258 586338 -5226 586894
rect -5846 550894 -5226 586338
rect -5846 550338 -5814 550894
rect -5258 550338 -5226 550894
rect -5846 514894 -5226 550338
rect -5846 514338 -5814 514894
rect -5258 514338 -5226 514894
rect -5846 478894 -5226 514338
rect -5846 478338 -5814 478894
rect -5258 478338 -5226 478894
rect -5846 442894 -5226 478338
rect -5846 442338 -5814 442894
rect -5258 442338 -5226 442894
rect -5846 406894 -5226 442338
rect -5846 406338 -5814 406894
rect -5258 406338 -5226 406894
rect -5846 370894 -5226 406338
rect -5846 370338 -5814 370894
rect -5258 370338 -5226 370894
rect -5846 334894 -5226 370338
rect -5846 334338 -5814 334894
rect -5258 334338 -5226 334894
rect -5846 298894 -5226 334338
rect -5846 298338 -5814 298894
rect -5258 298338 -5226 298894
rect -5846 262894 -5226 298338
rect -5846 262338 -5814 262894
rect -5258 262338 -5226 262894
rect -5846 226894 -5226 262338
rect -5846 226338 -5814 226894
rect -5258 226338 -5226 226894
rect -5846 190894 -5226 226338
rect -5846 190338 -5814 190894
rect -5258 190338 -5226 190894
rect -5846 154894 -5226 190338
rect -5846 154338 -5814 154894
rect -5258 154338 -5226 154894
rect -5846 118894 -5226 154338
rect -5846 118338 -5814 118894
rect -5258 118338 -5226 118894
rect -5846 82894 -5226 118338
rect -5846 82338 -5814 82894
rect -5258 82338 -5226 82894
rect -5846 46894 -5226 82338
rect -5846 46338 -5814 46894
rect -5258 46338 -5226 46894
rect -5846 10894 -5226 46338
rect -5846 10338 -5814 10894
rect -5258 10338 -5226 10894
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 673174 -4266 707162
rect -4886 672618 -4854 673174
rect -4298 672618 -4266 673174
rect -4886 637174 -4266 672618
rect -4886 636618 -4854 637174
rect -4298 636618 -4266 637174
rect -4886 601174 -4266 636618
rect -4886 600618 -4854 601174
rect -4298 600618 -4266 601174
rect -4886 565174 -4266 600618
rect -4886 564618 -4854 565174
rect -4298 564618 -4266 565174
rect -4886 529174 -4266 564618
rect -4886 528618 -4854 529174
rect -4298 528618 -4266 529174
rect -4886 493174 -4266 528618
rect -4886 492618 -4854 493174
rect -4298 492618 -4266 493174
rect -4886 457174 -4266 492618
rect -4886 456618 -4854 457174
rect -4298 456618 -4266 457174
rect -4886 421174 -4266 456618
rect -4886 420618 -4854 421174
rect -4298 420618 -4266 421174
rect -4886 385174 -4266 420618
rect -4886 384618 -4854 385174
rect -4298 384618 -4266 385174
rect -4886 349174 -4266 384618
rect -4886 348618 -4854 349174
rect -4298 348618 -4266 349174
rect -4886 313174 -4266 348618
rect -4886 312618 -4854 313174
rect -4298 312618 -4266 313174
rect -4886 277174 -4266 312618
rect -4886 276618 -4854 277174
rect -4298 276618 -4266 277174
rect -4886 241174 -4266 276618
rect -4886 240618 -4854 241174
rect -4298 240618 -4266 241174
rect -4886 205174 -4266 240618
rect -4886 204618 -4854 205174
rect -4298 204618 -4266 205174
rect -4886 169174 -4266 204618
rect -4886 168618 -4854 169174
rect -4298 168618 -4266 169174
rect -4886 133174 -4266 168618
rect -4886 132618 -4854 133174
rect -4298 132618 -4266 133174
rect -4886 97174 -4266 132618
rect -4886 96618 -4854 97174
rect -4298 96618 -4266 97174
rect -4886 61174 -4266 96618
rect -4886 60618 -4854 61174
rect -4298 60618 -4266 61174
rect -4886 25174 -4266 60618
rect -4886 24618 -4854 25174
rect -4298 24618 -4266 25174
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706202 5546 706758
rect 6102 706202 6134 706758
rect -3926 690618 -3894 691174
rect -3338 690618 -3306 691174
rect -3926 655174 -3306 690618
rect -3926 654618 -3894 655174
rect -3338 654618 -3306 655174
rect -3926 619174 -3306 654618
rect -3926 618618 -3894 619174
rect -3338 618618 -3306 619174
rect -3926 583174 -3306 618618
rect -3926 582618 -3894 583174
rect -3338 582618 -3306 583174
rect -3926 547174 -3306 582618
rect -3926 546618 -3894 547174
rect -3338 546618 -3306 547174
rect -3926 511174 -3306 546618
rect -3926 510618 -3894 511174
rect -3338 510618 -3306 511174
rect -3926 475174 -3306 510618
rect -3926 474618 -3894 475174
rect -3338 474618 -3306 475174
rect -3926 439174 -3306 474618
rect -3926 438618 -3894 439174
rect -3338 438618 -3306 439174
rect -3926 403174 -3306 438618
rect -3926 402618 -3894 403174
rect -3338 402618 -3306 403174
rect -3926 367174 -3306 402618
rect -3926 366618 -3894 367174
rect -3338 366618 -3306 367174
rect -3926 331174 -3306 366618
rect -3926 330618 -3894 331174
rect -3338 330618 -3306 331174
rect -3926 295174 -3306 330618
rect -3926 294618 -3894 295174
rect -3338 294618 -3306 295174
rect -3926 259174 -3306 294618
rect -3926 258618 -3894 259174
rect -3338 258618 -3306 259174
rect -3926 223174 -3306 258618
rect -3926 222618 -3894 223174
rect -3338 222618 -3306 223174
rect -3926 187174 -3306 222618
rect -3926 186618 -3894 187174
rect -3338 186618 -3306 187174
rect -3926 151174 -3306 186618
rect -3926 150618 -3894 151174
rect -3338 150618 -3306 151174
rect -3926 115174 -3306 150618
rect -3926 114618 -3894 115174
rect -3338 114618 -3306 115174
rect -3926 79174 -3306 114618
rect -3926 78618 -3894 79174
rect -3338 78618 -3306 79174
rect -3926 43174 -3306 78618
rect -3926 42618 -3894 43174
rect -3338 42618 -3306 43174
rect -3926 7174 -3306 42618
rect -3926 6618 -3894 7174
rect -3338 6618 -3306 7174
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 669454 -2346 705242
rect -2966 668898 -2934 669454
rect -2378 668898 -2346 669454
rect -2966 633454 -2346 668898
rect -2966 632898 -2934 633454
rect -2378 632898 -2346 633454
rect -2966 597454 -2346 632898
rect -2966 596898 -2934 597454
rect -2378 596898 -2346 597454
rect -2966 561454 -2346 596898
rect -2966 560898 -2934 561454
rect -2378 560898 -2346 561454
rect -2966 525454 -2346 560898
rect -2966 524898 -2934 525454
rect -2378 524898 -2346 525454
rect -2966 489454 -2346 524898
rect -2966 488898 -2934 489454
rect -2378 488898 -2346 489454
rect -2966 453454 -2346 488898
rect -2966 452898 -2934 453454
rect -2378 452898 -2346 453454
rect -2966 417454 -2346 452898
rect -2966 416898 -2934 417454
rect -2378 416898 -2346 417454
rect -2966 381454 -2346 416898
rect -2966 380898 -2934 381454
rect -2378 380898 -2346 381454
rect -2966 345454 -2346 380898
rect -2966 344898 -2934 345454
rect -2378 344898 -2346 345454
rect -2966 309454 -2346 344898
rect -2966 308898 -2934 309454
rect -2378 308898 -2346 309454
rect -2966 273454 -2346 308898
rect -2966 272898 -2934 273454
rect -2378 272898 -2346 273454
rect -2966 237454 -2346 272898
rect -2966 236898 -2934 237454
rect -2378 236898 -2346 237454
rect -2966 201454 -2346 236898
rect -2966 200898 -2934 201454
rect -2378 200898 -2346 201454
rect -2966 165454 -2346 200898
rect -2966 164898 -2934 165454
rect -2378 164898 -2346 165454
rect -2966 129454 -2346 164898
rect -2966 128898 -2934 129454
rect -2378 128898 -2346 129454
rect -2966 93454 -2346 128898
rect -2966 92898 -2934 93454
rect -2378 92898 -2346 93454
rect -2966 57454 -2346 92898
rect -2966 56898 -2934 57454
rect -2378 56898 -2346 57454
rect -2966 21454 -2346 56898
rect -2966 20898 -2934 21454
rect -2378 20898 -2346 21454
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 687454 -1386 704282
rect -2006 686898 -1974 687454
rect -1418 686898 -1386 687454
rect -2006 651454 -1386 686898
rect -2006 650898 -1974 651454
rect -1418 650898 -1386 651454
rect -2006 615454 -1386 650898
rect -2006 614898 -1974 615454
rect -1418 614898 -1386 615454
rect -2006 579454 -1386 614898
rect -2006 578898 -1974 579454
rect -1418 578898 -1386 579454
rect -2006 543454 -1386 578898
rect -2006 542898 -1974 543454
rect -1418 542898 -1386 543454
rect -2006 507454 -1386 542898
rect -2006 506898 -1974 507454
rect -1418 506898 -1386 507454
rect -2006 471454 -1386 506898
rect -2006 470898 -1974 471454
rect -1418 470898 -1386 471454
rect -2006 435454 -1386 470898
rect -2006 434898 -1974 435454
rect -1418 434898 -1386 435454
rect -2006 399454 -1386 434898
rect -2006 398898 -1974 399454
rect -1418 398898 -1386 399454
rect -2006 363454 -1386 398898
rect -2006 362898 -1974 363454
rect -1418 362898 -1386 363454
rect -2006 327454 -1386 362898
rect -2006 326898 -1974 327454
rect -1418 326898 -1386 327454
rect -2006 291454 -1386 326898
rect -2006 290898 -1974 291454
rect -1418 290898 -1386 291454
rect -2006 255454 -1386 290898
rect -2006 254898 -1974 255454
rect -1418 254898 -1386 255454
rect -2006 219454 -1386 254898
rect -2006 218898 -1974 219454
rect -1418 218898 -1386 219454
rect -2006 183454 -1386 218898
rect -2006 182898 -1974 183454
rect -1418 182898 -1386 183454
rect -2006 147454 -1386 182898
rect -2006 146898 -1974 147454
rect -1418 146898 -1386 147454
rect -2006 111454 -1386 146898
rect -2006 110898 -1974 111454
rect -1418 110898 -1386 111454
rect -2006 75454 -1386 110898
rect -2006 74898 -1974 75454
rect -1418 74898 -1386 75454
rect -2006 39454 -1386 74898
rect -2006 38898 -1974 39454
rect -1418 38898 -1386 39454
rect -2006 3454 -1386 38898
rect -2006 2898 -1974 3454
rect -1418 2898 -1386 3454
rect -2006 -346 -1386 2898
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704282 1826 704838
rect 2382 704282 2414 704838
rect 1794 687454 2414 704282
rect 1794 686898 1826 687454
rect 2382 686898 2414 687454
rect 1794 651454 2414 686898
rect 1794 650898 1826 651454
rect 2382 650898 2414 651454
rect 1794 615454 2414 650898
rect 1794 614898 1826 615454
rect 2382 614898 2414 615454
rect 1794 579454 2414 614898
rect 1794 578898 1826 579454
rect 2382 578898 2414 579454
rect 1794 543454 2414 578898
rect 1794 542898 1826 543454
rect 2382 542898 2414 543454
rect 1794 507454 2414 542898
rect 1794 506898 1826 507454
rect 2382 506898 2414 507454
rect 1794 471454 2414 506898
rect 1794 470898 1826 471454
rect 2382 470898 2414 471454
rect 1794 435454 2414 470898
rect 1794 434898 1826 435454
rect 2382 434898 2414 435454
rect 1794 399454 2414 434898
rect 1794 398898 1826 399454
rect 2382 398898 2414 399454
rect 1794 363454 2414 398898
rect 1794 362898 1826 363454
rect 2382 362898 2414 363454
rect 1794 327454 2414 362898
rect 1794 326898 1826 327454
rect 2382 326898 2414 327454
rect 1794 291454 2414 326898
rect 1794 290898 1826 291454
rect 2382 290898 2414 291454
rect 1794 255454 2414 290898
rect 1794 254898 1826 255454
rect 2382 254898 2414 255454
rect 1794 219454 2414 254898
rect 1794 218898 1826 219454
rect 2382 218898 2414 219454
rect 1794 183454 2414 218898
rect 1794 182898 1826 183454
rect 2382 182898 2414 183454
rect 1794 147454 2414 182898
rect 1794 146898 1826 147454
rect 2382 146898 2414 147454
rect 1794 111454 2414 146898
rect 1794 110898 1826 111454
rect 2382 110898 2414 111454
rect 1794 75454 2414 110898
rect 1794 74898 1826 75454
rect 2382 74898 2414 75454
rect 1794 39454 2414 74898
rect 1794 38898 1826 39454
rect 2382 38898 2414 39454
rect 1794 3454 2414 38898
rect 1794 2898 1826 3454
rect 2382 2898 2414 3454
rect 1794 -346 2414 2898
rect 1794 -902 1826 -346
rect 2382 -902 2414 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690618 5546 691174
rect 6102 690618 6134 691174
rect 5514 655174 6134 690618
rect 5514 654618 5546 655174
rect 6102 654618 6134 655174
rect 5514 619174 6134 654618
rect 5514 618618 5546 619174
rect 6102 618618 6134 619174
rect 5514 583174 6134 618618
rect 5514 582618 5546 583174
rect 6102 582618 6134 583174
rect 5514 547174 6134 582618
rect 5514 546618 5546 547174
rect 6102 546618 6134 547174
rect 5514 511174 6134 546618
rect 5514 510618 5546 511174
rect 6102 510618 6134 511174
rect 5514 475174 6134 510618
rect 5514 474618 5546 475174
rect 6102 474618 6134 475174
rect 5514 439174 6134 474618
rect 5514 438618 5546 439174
rect 6102 438618 6134 439174
rect 5514 403174 6134 438618
rect 5514 402618 5546 403174
rect 6102 402618 6134 403174
rect 5514 367174 6134 402618
rect 5514 366618 5546 367174
rect 6102 366618 6134 367174
rect 5514 331174 6134 366618
rect 5514 330618 5546 331174
rect 6102 330618 6134 331174
rect 5514 295174 6134 330618
rect 5514 294618 5546 295174
rect 6102 294618 6134 295174
rect 5514 259174 6134 294618
rect 5514 258618 5546 259174
rect 6102 258618 6134 259174
rect 5514 223174 6134 258618
rect 5514 222618 5546 223174
rect 6102 222618 6134 223174
rect 5514 187174 6134 222618
rect 5514 186618 5546 187174
rect 6102 186618 6134 187174
rect 5514 151174 6134 186618
rect 5514 150618 5546 151174
rect 6102 150618 6134 151174
rect 5514 115174 6134 150618
rect 5514 114618 5546 115174
rect 6102 114618 6134 115174
rect 5514 79174 6134 114618
rect 5514 78618 5546 79174
rect 6102 78618 6134 79174
rect 5514 43174 6134 78618
rect 5514 42618 5546 43174
rect 6102 42618 6134 43174
rect 5514 7174 6134 42618
rect 5514 6618 5546 7174
rect 6102 6618 6134 7174
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2822 5546 -2266
rect 6102 -2822 6134 -2266
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694338 9266 694894
rect 9822 694338 9854 694894
rect 9234 658894 9854 694338
rect 9234 658338 9266 658894
rect 9822 658338 9854 658894
rect 9234 622894 9854 658338
rect 9234 622338 9266 622894
rect 9822 622338 9854 622894
rect 9234 586894 9854 622338
rect 9234 586338 9266 586894
rect 9822 586338 9854 586894
rect 9234 550894 9854 586338
rect 9234 550338 9266 550894
rect 9822 550338 9854 550894
rect 9234 514894 9854 550338
rect 9234 514338 9266 514894
rect 9822 514338 9854 514894
rect 9234 478894 9854 514338
rect 9234 478338 9266 478894
rect 9822 478338 9854 478894
rect 9234 442894 9854 478338
rect 9234 442338 9266 442894
rect 9822 442338 9854 442894
rect 9234 406894 9854 442338
rect 9234 406338 9266 406894
rect 9822 406338 9854 406894
rect 9234 370894 9854 406338
rect 9234 370338 9266 370894
rect 9822 370338 9854 370894
rect 9234 334894 9854 370338
rect 9234 334338 9266 334894
rect 9822 334338 9854 334894
rect 9234 298894 9854 334338
rect 9234 298338 9266 298894
rect 9822 298338 9854 298894
rect 9234 262894 9854 298338
rect 9234 262338 9266 262894
rect 9822 262338 9854 262894
rect 9234 226894 9854 262338
rect 9234 226338 9266 226894
rect 9822 226338 9854 226894
rect 9234 190894 9854 226338
rect 9234 190338 9266 190894
rect 9822 190338 9854 190894
rect 9234 154894 9854 190338
rect 9234 154338 9266 154894
rect 9822 154338 9854 154894
rect 9234 118894 9854 154338
rect 9234 118338 9266 118894
rect 9822 118338 9854 118894
rect 9234 82894 9854 118338
rect 9234 82338 9266 82894
rect 9822 82338 9854 82894
rect 9234 46894 9854 82338
rect 9234 46338 9266 46894
rect 9822 46338 9854 46894
rect 9234 10894 9854 46338
rect 9234 10338 9266 10894
rect 9822 10338 9854 10894
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4742 9266 -4186
rect 9822 -4742 9854 -4186
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711002 30986 711558
rect 31542 711002 31574 711558
rect 27234 709638 27854 709670
rect 27234 709082 27266 709638
rect 27822 709082 27854 709638
rect 23514 707718 24134 707750
rect 23514 707162 23546 707718
rect 24102 707162 24134 707718
rect 12954 698058 12986 698614
rect 13542 698058 13574 698614
rect 12954 662614 13574 698058
rect 12954 662058 12986 662614
rect 13542 662058 13574 662614
rect 12954 626614 13574 662058
rect 12954 626058 12986 626614
rect 13542 626058 13574 626614
rect 12954 590614 13574 626058
rect 12954 590058 12986 590614
rect 13542 590058 13574 590614
rect 12954 554614 13574 590058
rect 12954 554058 12986 554614
rect 13542 554058 13574 554614
rect 12954 518614 13574 554058
rect 12954 518058 12986 518614
rect 13542 518058 13574 518614
rect 12954 482614 13574 518058
rect 12954 482058 12986 482614
rect 13542 482058 13574 482614
rect 12954 446614 13574 482058
rect 12954 446058 12986 446614
rect 13542 446058 13574 446614
rect 12954 410614 13574 446058
rect 12954 410058 12986 410614
rect 13542 410058 13574 410614
rect 12954 374614 13574 410058
rect 12954 374058 12986 374614
rect 13542 374058 13574 374614
rect 12954 338614 13574 374058
rect 12954 338058 12986 338614
rect 13542 338058 13574 338614
rect 12954 302614 13574 338058
rect 12954 302058 12986 302614
rect 13542 302058 13574 302614
rect 12954 266614 13574 302058
rect 12954 266058 12986 266614
rect 13542 266058 13574 266614
rect 12954 230614 13574 266058
rect 12954 230058 12986 230614
rect 13542 230058 13574 230614
rect 12954 194614 13574 230058
rect 12954 194058 12986 194614
rect 13542 194058 13574 194614
rect 12954 158614 13574 194058
rect 12954 158058 12986 158614
rect 13542 158058 13574 158614
rect 12954 122614 13574 158058
rect 12954 122058 12986 122614
rect 13542 122058 13574 122614
rect 12954 86614 13574 122058
rect 12954 86058 12986 86614
rect 13542 86058 13574 86614
rect 12954 50614 13574 86058
rect 12954 50058 12986 50614
rect 13542 50058 13574 50614
rect 12954 14614 13574 50058
rect 12954 14058 12986 14614
rect 13542 14058 13574 14614
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705242 19826 705798
rect 20382 705242 20414 705798
rect 19794 669454 20414 705242
rect 19794 668898 19826 669454
rect 20382 668898 20414 669454
rect 19794 633454 20414 668898
rect 19794 632898 19826 633454
rect 20382 632898 20414 633454
rect 19794 597454 20414 632898
rect 19794 596898 19826 597454
rect 20382 596898 20414 597454
rect 19794 561454 20414 596898
rect 19794 560898 19826 561454
rect 20382 560898 20414 561454
rect 19794 525454 20414 560898
rect 19794 524898 19826 525454
rect 20382 524898 20414 525454
rect 19794 489454 20414 524898
rect 19794 488898 19826 489454
rect 20382 488898 20414 489454
rect 19794 453454 20414 488898
rect 19794 452898 19826 453454
rect 20382 452898 20414 453454
rect 19794 417454 20414 452898
rect 19794 416898 19826 417454
rect 20382 416898 20414 417454
rect 19794 381454 20414 416898
rect 19794 380898 19826 381454
rect 20382 380898 20414 381454
rect 19794 345454 20414 380898
rect 19794 344898 19826 345454
rect 20382 344898 20414 345454
rect 19794 309454 20414 344898
rect 19794 308898 19826 309454
rect 20382 308898 20414 309454
rect 19794 273454 20414 308898
rect 19794 272898 19826 273454
rect 20382 272898 20414 273454
rect 19794 237454 20414 272898
rect 19794 236898 19826 237454
rect 20382 236898 20414 237454
rect 19794 201454 20414 236898
rect 19794 200898 19826 201454
rect 20382 200898 20414 201454
rect 19794 165454 20414 200898
rect 19794 164898 19826 165454
rect 20382 164898 20414 165454
rect 19794 129454 20414 164898
rect 19794 128898 19826 129454
rect 20382 128898 20414 129454
rect 19794 93454 20414 128898
rect 19794 92898 19826 93454
rect 20382 92898 20414 93454
rect 19794 57454 20414 92898
rect 19794 56898 19826 57454
rect 20382 56898 20414 57454
rect 19794 21454 20414 56898
rect 19794 20898 19826 21454
rect 20382 20898 20414 21454
rect 19794 -1306 20414 20898
rect 19794 -1862 19826 -1306
rect 20382 -1862 20414 -1306
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672618 23546 673174
rect 24102 672618 24134 673174
rect 23514 637174 24134 672618
rect 23514 636618 23546 637174
rect 24102 636618 24134 637174
rect 23514 601174 24134 636618
rect 23514 600618 23546 601174
rect 24102 600618 24134 601174
rect 23514 565174 24134 600618
rect 23514 564618 23546 565174
rect 24102 564618 24134 565174
rect 23514 529174 24134 564618
rect 23514 528618 23546 529174
rect 24102 528618 24134 529174
rect 23514 493174 24134 528618
rect 23514 492618 23546 493174
rect 24102 492618 24134 493174
rect 23514 457174 24134 492618
rect 23514 456618 23546 457174
rect 24102 456618 24134 457174
rect 23514 421174 24134 456618
rect 23514 420618 23546 421174
rect 24102 420618 24134 421174
rect 23514 385174 24134 420618
rect 23514 384618 23546 385174
rect 24102 384618 24134 385174
rect 23514 349174 24134 384618
rect 23514 348618 23546 349174
rect 24102 348618 24134 349174
rect 23514 313174 24134 348618
rect 23514 312618 23546 313174
rect 24102 312618 24134 313174
rect 23514 277174 24134 312618
rect 23514 276618 23546 277174
rect 24102 276618 24134 277174
rect 23514 241174 24134 276618
rect 23514 240618 23546 241174
rect 24102 240618 24134 241174
rect 23514 205174 24134 240618
rect 23514 204618 23546 205174
rect 24102 204618 24134 205174
rect 23514 169174 24134 204618
rect 23514 168618 23546 169174
rect 24102 168618 24134 169174
rect 23514 133174 24134 168618
rect 23514 132618 23546 133174
rect 24102 132618 24134 133174
rect 23514 97174 24134 132618
rect 23514 96618 23546 97174
rect 24102 96618 24134 97174
rect 23514 61174 24134 96618
rect 23514 60618 23546 61174
rect 24102 60618 24134 61174
rect 23514 25174 24134 60618
rect 23514 24618 23546 25174
rect 24102 24618 24134 25174
rect 23514 -3226 24134 24618
rect 23514 -3782 23546 -3226
rect 24102 -3782 24134 -3226
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676338 27266 676894
rect 27822 676338 27854 676894
rect 27234 640894 27854 676338
rect 27234 640338 27266 640894
rect 27822 640338 27854 640894
rect 27234 604894 27854 640338
rect 27234 604338 27266 604894
rect 27822 604338 27854 604894
rect 27234 568894 27854 604338
rect 27234 568338 27266 568894
rect 27822 568338 27854 568894
rect 27234 532894 27854 568338
rect 27234 532338 27266 532894
rect 27822 532338 27854 532894
rect 27234 496894 27854 532338
rect 27234 496338 27266 496894
rect 27822 496338 27854 496894
rect 27234 460894 27854 496338
rect 27234 460338 27266 460894
rect 27822 460338 27854 460894
rect 27234 424894 27854 460338
rect 27234 424338 27266 424894
rect 27822 424338 27854 424894
rect 27234 388894 27854 424338
rect 27234 388338 27266 388894
rect 27822 388338 27854 388894
rect 27234 352894 27854 388338
rect 27234 352338 27266 352894
rect 27822 352338 27854 352894
rect 27234 316894 27854 352338
rect 27234 316338 27266 316894
rect 27822 316338 27854 316894
rect 27234 280894 27854 316338
rect 27234 280338 27266 280894
rect 27822 280338 27854 280894
rect 27234 244894 27854 280338
rect 27234 244338 27266 244894
rect 27822 244338 27854 244894
rect 27234 208894 27854 244338
rect 27234 208338 27266 208894
rect 27822 208338 27854 208894
rect 27234 172894 27854 208338
rect 27234 172338 27266 172894
rect 27822 172338 27854 172894
rect 27234 136894 27854 172338
rect 27234 136338 27266 136894
rect 27822 136338 27854 136894
rect 27234 100894 27854 136338
rect 27234 100338 27266 100894
rect 27822 100338 27854 100894
rect 27234 64894 27854 100338
rect 27234 64338 27266 64894
rect 27822 64338 27854 64894
rect 27234 28894 27854 64338
rect 27234 28338 27266 28894
rect 27822 28338 27854 28894
rect 27234 -5146 27854 28338
rect 27234 -5702 27266 -5146
rect 27822 -5702 27854 -5146
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710042 48986 710598
rect 49542 710042 49574 710598
rect 45234 708678 45854 709670
rect 45234 708122 45266 708678
rect 45822 708122 45854 708678
rect 41514 706758 42134 707750
rect 41514 706202 41546 706758
rect 42102 706202 42134 706758
rect 30954 680058 30986 680614
rect 31542 680058 31574 680614
rect 30954 644614 31574 680058
rect 30954 644058 30986 644614
rect 31542 644058 31574 644614
rect 30954 608614 31574 644058
rect 30954 608058 30986 608614
rect 31542 608058 31574 608614
rect 30954 572614 31574 608058
rect 30954 572058 30986 572614
rect 31542 572058 31574 572614
rect 30954 536614 31574 572058
rect 30954 536058 30986 536614
rect 31542 536058 31574 536614
rect 30954 500614 31574 536058
rect 30954 500058 30986 500614
rect 31542 500058 31574 500614
rect 30954 464614 31574 500058
rect 30954 464058 30986 464614
rect 31542 464058 31574 464614
rect 30954 428614 31574 464058
rect 30954 428058 30986 428614
rect 31542 428058 31574 428614
rect 30954 392614 31574 428058
rect 30954 392058 30986 392614
rect 31542 392058 31574 392614
rect 30954 356614 31574 392058
rect 30954 356058 30986 356614
rect 31542 356058 31574 356614
rect 30954 320614 31574 356058
rect 30954 320058 30986 320614
rect 31542 320058 31574 320614
rect 30954 284614 31574 320058
rect 30954 284058 30986 284614
rect 31542 284058 31574 284614
rect 30954 248614 31574 284058
rect 30954 248058 30986 248614
rect 31542 248058 31574 248614
rect 30954 212614 31574 248058
rect 30954 212058 30986 212614
rect 31542 212058 31574 212614
rect 30954 176614 31574 212058
rect 30954 176058 30986 176614
rect 31542 176058 31574 176614
rect 30954 140614 31574 176058
rect 30954 140058 30986 140614
rect 31542 140058 31574 140614
rect 30954 104614 31574 140058
rect 30954 104058 30986 104614
rect 31542 104058 31574 104614
rect 30954 68614 31574 104058
rect 30954 68058 30986 68614
rect 31542 68058 31574 68614
rect 30954 32614 31574 68058
rect 30954 32058 30986 32614
rect 31542 32058 31574 32614
rect 12954 -6662 12986 -6106
rect 13542 -6662 13574 -6106
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704282 37826 704838
rect 38382 704282 38414 704838
rect 37794 687454 38414 704282
rect 37794 686898 37826 687454
rect 38382 686898 38414 687454
rect 37794 651454 38414 686898
rect 37794 650898 37826 651454
rect 38382 650898 38414 651454
rect 37794 615454 38414 650898
rect 37794 614898 37826 615454
rect 38382 614898 38414 615454
rect 37794 579454 38414 614898
rect 37794 578898 37826 579454
rect 38382 578898 38414 579454
rect 37794 543454 38414 578898
rect 37794 542898 37826 543454
rect 38382 542898 38414 543454
rect 37794 507454 38414 542898
rect 37794 506898 37826 507454
rect 38382 506898 38414 507454
rect 37794 471454 38414 506898
rect 37794 470898 37826 471454
rect 38382 470898 38414 471454
rect 37794 435454 38414 470898
rect 37794 434898 37826 435454
rect 38382 434898 38414 435454
rect 37794 399454 38414 434898
rect 37794 398898 37826 399454
rect 38382 398898 38414 399454
rect 37794 363454 38414 398898
rect 37794 362898 37826 363454
rect 38382 362898 38414 363454
rect 37794 327454 38414 362898
rect 37794 326898 37826 327454
rect 38382 326898 38414 327454
rect 37794 291454 38414 326898
rect 37794 290898 37826 291454
rect 38382 290898 38414 291454
rect 37794 255454 38414 290898
rect 37794 254898 37826 255454
rect 38382 254898 38414 255454
rect 37794 219454 38414 254898
rect 37794 218898 37826 219454
rect 38382 218898 38414 219454
rect 37794 183454 38414 218898
rect 37794 182898 37826 183454
rect 38382 182898 38414 183454
rect 37794 147454 38414 182898
rect 37794 146898 37826 147454
rect 38382 146898 38414 147454
rect 37794 111454 38414 146898
rect 37794 110898 37826 111454
rect 38382 110898 38414 111454
rect 37794 75454 38414 110898
rect 37794 74898 37826 75454
rect 38382 74898 38414 75454
rect 37794 39454 38414 74898
rect 37794 38898 37826 39454
rect 38382 38898 38414 39454
rect 37794 3454 38414 38898
rect 37794 2898 37826 3454
rect 38382 2898 38414 3454
rect 37794 -346 38414 2898
rect 37794 -902 37826 -346
rect 38382 -902 38414 -346
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690618 41546 691174
rect 42102 690618 42134 691174
rect 41514 655174 42134 690618
rect 41514 654618 41546 655174
rect 42102 654618 42134 655174
rect 41514 619174 42134 654618
rect 41514 618618 41546 619174
rect 42102 618618 42134 619174
rect 41514 583174 42134 618618
rect 41514 582618 41546 583174
rect 42102 582618 42134 583174
rect 41514 547174 42134 582618
rect 41514 546618 41546 547174
rect 42102 546618 42134 547174
rect 41514 511174 42134 546618
rect 41514 510618 41546 511174
rect 42102 510618 42134 511174
rect 41514 475174 42134 510618
rect 41514 474618 41546 475174
rect 42102 474618 42134 475174
rect 41514 439174 42134 474618
rect 41514 438618 41546 439174
rect 42102 438618 42134 439174
rect 41514 403174 42134 438618
rect 41514 402618 41546 403174
rect 42102 402618 42134 403174
rect 41514 367174 42134 402618
rect 41514 366618 41546 367174
rect 42102 366618 42134 367174
rect 41514 331174 42134 366618
rect 41514 330618 41546 331174
rect 42102 330618 42134 331174
rect 41514 295174 42134 330618
rect 41514 294618 41546 295174
rect 42102 294618 42134 295174
rect 41514 259174 42134 294618
rect 41514 258618 41546 259174
rect 42102 258618 42134 259174
rect 41514 223174 42134 258618
rect 41514 222618 41546 223174
rect 42102 222618 42134 223174
rect 41514 187174 42134 222618
rect 41514 186618 41546 187174
rect 42102 186618 42134 187174
rect 41514 151174 42134 186618
rect 41514 150618 41546 151174
rect 42102 150618 42134 151174
rect 41514 115174 42134 150618
rect 41514 114618 41546 115174
rect 42102 114618 42134 115174
rect 41514 79174 42134 114618
rect 41514 78618 41546 79174
rect 42102 78618 42134 79174
rect 41514 43174 42134 78618
rect 41514 42618 41546 43174
rect 42102 42618 42134 43174
rect 41514 7174 42134 42618
rect 41514 6618 41546 7174
rect 42102 6618 42134 7174
rect 41514 -2266 42134 6618
rect 41514 -2822 41546 -2266
rect 42102 -2822 42134 -2266
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694338 45266 694894
rect 45822 694338 45854 694894
rect 45234 658894 45854 694338
rect 45234 658338 45266 658894
rect 45822 658338 45854 658894
rect 45234 622894 45854 658338
rect 45234 622338 45266 622894
rect 45822 622338 45854 622894
rect 45234 586894 45854 622338
rect 45234 586338 45266 586894
rect 45822 586338 45854 586894
rect 45234 550894 45854 586338
rect 45234 550338 45266 550894
rect 45822 550338 45854 550894
rect 45234 514894 45854 550338
rect 45234 514338 45266 514894
rect 45822 514338 45854 514894
rect 45234 478894 45854 514338
rect 45234 478338 45266 478894
rect 45822 478338 45854 478894
rect 45234 442894 45854 478338
rect 45234 442338 45266 442894
rect 45822 442338 45854 442894
rect 45234 406894 45854 442338
rect 45234 406338 45266 406894
rect 45822 406338 45854 406894
rect 45234 370894 45854 406338
rect 45234 370338 45266 370894
rect 45822 370338 45854 370894
rect 45234 334894 45854 370338
rect 45234 334338 45266 334894
rect 45822 334338 45854 334894
rect 45234 298894 45854 334338
rect 45234 298338 45266 298894
rect 45822 298338 45854 298894
rect 45234 262894 45854 298338
rect 45234 262338 45266 262894
rect 45822 262338 45854 262894
rect 45234 226894 45854 262338
rect 45234 226338 45266 226894
rect 45822 226338 45854 226894
rect 45234 190894 45854 226338
rect 45234 190338 45266 190894
rect 45822 190338 45854 190894
rect 45234 154894 45854 190338
rect 45234 154338 45266 154894
rect 45822 154338 45854 154894
rect 45234 118894 45854 154338
rect 45234 118338 45266 118894
rect 45822 118338 45854 118894
rect 45234 82894 45854 118338
rect 45234 82338 45266 82894
rect 45822 82338 45854 82894
rect 45234 46894 45854 82338
rect 45234 46338 45266 46894
rect 45822 46338 45854 46894
rect 45234 10894 45854 46338
rect 45234 10338 45266 10894
rect 45822 10338 45854 10894
rect 45234 -4186 45854 10338
rect 45234 -4742 45266 -4186
rect 45822 -4742 45854 -4186
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711002 66986 711558
rect 67542 711002 67574 711558
rect 63234 709638 63854 709670
rect 63234 709082 63266 709638
rect 63822 709082 63854 709638
rect 59514 707718 60134 707750
rect 59514 707162 59546 707718
rect 60102 707162 60134 707718
rect 48954 698058 48986 698614
rect 49542 698058 49574 698614
rect 48954 662614 49574 698058
rect 48954 662058 48986 662614
rect 49542 662058 49574 662614
rect 48954 626614 49574 662058
rect 48954 626058 48986 626614
rect 49542 626058 49574 626614
rect 48954 590614 49574 626058
rect 48954 590058 48986 590614
rect 49542 590058 49574 590614
rect 48954 554614 49574 590058
rect 48954 554058 48986 554614
rect 49542 554058 49574 554614
rect 48954 518614 49574 554058
rect 48954 518058 48986 518614
rect 49542 518058 49574 518614
rect 48954 482614 49574 518058
rect 48954 482058 48986 482614
rect 49542 482058 49574 482614
rect 48954 446614 49574 482058
rect 48954 446058 48986 446614
rect 49542 446058 49574 446614
rect 48954 410614 49574 446058
rect 48954 410058 48986 410614
rect 49542 410058 49574 410614
rect 48954 374614 49574 410058
rect 48954 374058 48986 374614
rect 49542 374058 49574 374614
rect 48954 338614 49574 374058
rect 48954 338058 48986 338614
rect 49542 338058 49574 338614
rect 48954 302614 49574 338058
rect 48954 302058 48986 302614
rect 49542 302058 49574 302614
rect 48954 266614 49574 302058
rect 48954 266058 48986 266614
rect 49542 266058 49574 266614
rect 48954 230614 49574 266058
rect 48954 230058 48986 230614
rect 49542 230058 49574 230614
rect 48954 194614 49574 230058
rect 48954 194058 48986 194614
rect 49542 194058 49574 194614
rect 48954 158614 49574 194058
rect 48954 158058 48986 158614
rect 49542 158058 49574 158614
rect 48954 122614 49574 158058
rect 48954 122058 48986 122614
rect 49542 122058 49574 122614
rect 48954 86614 49574 122058
rect 48954 86058 48986 86614
rect 49542 86058 49574 86614
rect 48954 50614 49574 86058
rect 48954 50058 48986 50614
rect 49542 50058 49574 50614
rect 48954 14614 49574 50058
rect 48954 14058 48986 14614
rect 49542 14058 49574 14614
rect 30954 -7622 30986 -7066
rect 31542 -7622 31574 -7066
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705242 55826 705798
rect 56382 705242 56414 705798
rect 55794 669454 56414 705242
rect 55794 668898 55826 669454
rect 56382 668898 56414 669454
rect 55794 633454 56414 668898
rect 55794 632898 55826 633454
rect 56382 632898 56414 633454
rect 55794 597454 56414 632898
rect 55794 596898 55826 597454
rect 56382 596898 56414 597454
rect 55794 561454 56414 596898
rect 55794 560898 55826 561454
rect 56382 560898 56414 561454
rect 55794 525454 56414 560898
rect 55794 524898 55826 525454
rect 56382 524898 56414 525454
rect 55794 489454 56414 524898
rect 55794 488898 55826 489454
rect 56382 488898 56414 489454
rect 55794 453454 56414 488898
rect 55794 452898 55826 453454
rect 56382 452898 56414 453454
rect 55794 417454 56414 452898
rect 55794 416898 55826 417454
rect 56382 416898 56414 417454
rect 55794 381454 56414 416898
rect 55794 380898 55826 381454
rect 56382 380898 56414 381454
rect 55794 345454 56414 380898
rect 55794 344898 55826 345454
rect 56382 344898 56414 345454
rect 55794 309454 56414 344898
rect 55794 308898 55826 309454
rect 56382 308898 56414 309454
rect 55794 273454 56414 308898
rect 55794 272898 55826 273454
rect 56382 272898 56414 273454
rect 55794 237454 56414 272898
rect 55794 236898 55826 237454
rect 56382 236898 56414 237454
rect 55794 201454 56414 236898
rect 55794 200898 55826 201454
rect 56382 200898 56414 201454
rect 55794 165454 56414 200898
rect 55794 164898 55826 165454
rect 56382 164898 56414 165454
rect 55794 129454 56414 164898
rect 55794 128898 55826 129454
rect 56382 128898 56414 129454
rect 55794 93454 56414 128898
rect 55794 92898 55826 93454
rect 56382 92898 56414 93454
rect 55794 57454 56414 92898
rect 55794 56898 55826 57454
rect 56382 56898 56414 57454
rect 55794 21454 56414 56898
rect 55794 20898 55826 21454
rect 56382 20898 56414 21454
rect 55794 -1306 56414 20898
rect 55794 -1862 55826 -1306
rect 56382 -1862 56414 -1306
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672618 59546 673174
rect 60102 672618 60134 673174
rect 59514 637174 60134 672618
rect 59514 636618 59546 637174
rect 60102 636618 60134 637174
rect 59514 601174 60134 636618
rect 59514 600618 59546 601174
rect 60102 600618 60134 601174
rect 59514 565174 60134 600618
rect 59514 564618 59546 565174
rect 60102 564618 60134 565174
rect 59514 529174 60134 564618
rect 59514 528618 59546 529174
rect 60102 528618 60134 529174
rect 59514 493174 60134 528618
rect 59514 492618 59546 493174
rect 60102 492618 60134 493174
rect 59514 457174 60134 492618
rect 59514 456618 59546 457174
rect 60102 456618 60134 457174
rect 59514 421174 60134 456618
rect 59514 420618 59546 421174
rect 60102 420618 60134 421174
rect 59514 385174 60134 420618
rect 59514 384618 59546 385174
rect 60102 384618 60134 385174
rect 59514 349174 60134 384618
rect 59514 348618 59546 349174
rect 60102 348618 60134 349174
rect 59514 313174 60134 348618
rect 59514 312618 59546 313174
rect 60102 312618 60134 313174
rect 59514 277174 60134 312618
rect 59514 276618 59546 277174
rect 60102 276618 60134 277174
rect 59514 241174 60134 276618
rect 59514 240618 59546 241174
rect 60102 240618 60134 241174
rect 59514 205174 60134 240618
rect 59514 204618 59546 205174
rect 60102 204618 60134 205174
rect 59514 169174 60134 204618
rect 59514 168618 59546 169174
rect 60102 168618 60134 169174
rect 59514 133174 60134 168618
rect 59514 132618 59546 133174
rect 60102 132618 60134 133174
rect 59514 97174 60134 132618
rect 59514 96618 59546 97174
rect 60102 96618 60134 97174
rect 59514 61174 60134 96618
rect 59514 60618 59546 61174
rect 60102 60618 60134 61174
rect 59514 25174 60134 60618
rect 59514 24618 59546 25174
rect 60102 24618 60134 25174
rect 59514 -3226 60134 24618
rect 59514 -3782 59546 -3226
rect 60102 -3782 60134 -3226
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676338 63266 676894
rect 63822 676338 63854 676894
rect 63234 640894 63854 676338
rect 63234 640338 63266 640894
rect 63822 640338 63854 640894
rect 63234 604894 63854 640338
rect 63234 604338 63266 604894
rect 63822 604338 63854 604894
rect 63234 568894 63854 604338
rect 63234 568338 63266 568894
rect 63822 568338 63854 568894
rect 63234 532894 63854 568338
rect 63234 532338 63266 532894
rect 63822 532338 63854 532894
rect 63234 496894 63854 532338
rect 63234 496338 63266 496894
rect 63822 496338 63854 496894
rect 63234 460894 63854 496338
rect 63234 460338 63266 460894
rect 63822 460338 63854 460894
rect 63234 424894 63854 460338
rect 63234 424338 63266 424894
rect 63822 424338 63854 424894
rect 63234 388894 63854 424338
rect 63234 388338 63266 388894
rect 63822 388338 63854 388894
rect 63234 352894 63854 388338
rect 63234 352338 63266 352894
rect 63822 352338 63854 352894
rect 63234 316894 63854 352338
rect 63234 316338 63266 316894
rect 63822 316338 63854 316894
rect 63234 280894 63854 316338
rect 63234 280338 63266 280894
rect 63822 280338 63854 280894
rect 63234 244894 63854 280338
rect 63234 244338 63266 244894
rect 63822 244338 63854 244894
rect 63234 208894 63854 244338
rect 63234 208338 63266 208894
rect 63822 208338 63854 208894
rect 63234 172894 63854 208338
rect 63234 172338 63266 172894
rect 63822 172338 63854 172894
rect 63234 136894 63854 172338
rect 63234 136338 63266 136894
rect 63822 136338 63854 136894
rect 63234 100894 63854 136338
rect 63234 100338 63266 100894
rect 63822 100338 63854 100894
rect 63234 64894 63854 100338
rect 63234 64338 63266 64894
rect 63822 64338 63854 64894
rect 63234 28894 63854 64338
rect 63234 28338 63266 28894
rect 63822 28338 63854 28894
rect 63234 -5146 63854 28338
rect 63234 -5702 63266 -5146
rect 63822 -5702 63854 -5146
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710042 84986 710598
rect 85542 710042 85574 710598
rect 81234 708678 81854 709670
rect 81234 708122 81266 708678
rect 81822 708122 81854 708678
rect 77514 706758 78134 707750
rect 77514 706202 77546 706758
rect 78102 706202 78134 706758
rect 66954 680058 66986 680614
rect 67542 680058 67574 680614
rect 66954 644614 67574 680058
rect 66954 644058 66986 644614
rect 67542 644058 67574 644614
rect 66954 608614 67574 644058
rect 66954 608058 66986 608614
rect 67542 608058 67574 608614
rect 66954 572614 67574 608058
rect 66954 572058 66986 572614
rect 67542 572058 67574 572614
rect 66954 536614 67574 572058
rect 66954 536058 66986 536614
rect 67542 536058 67574 536614
rect 66954 500614 67574 536058
rect 66954 500058 66986 500614
rect 67542 500058 67574 500614
rect 66954 464614 67574 500058
rect 66954 464058 66986 464614
rect 67542 464058 67574 464614
rect 66954 428614 67574 464058
rect 66954 428058 66986 428614
rect 67542 428058 67574 428614
rect 66954 392614 67574 428058
rect 66954 392058 66986 392614
rect 67542 392058 67574 392614
rect 66954 356614 67574 392058
rect 66954 356058 66986 356614
rect 67542 356058 67574 356614
rect 66954 320614 67574 356058
rect 66954 320058 66986 320614
rect 67542 320058 67574 320614
rect 66954 284614 67574 320058
rect 66954 284058 66986 284614
rect 67542 284058 67574 284614
rect 66954 248614 67574 284058
rect 66954 248058 66986 248614
rect 67542 248058 67574 248614
rect 66954 212614 67574 248058
rect 66954 212058 66986 212614
rect 67542 212058 67574 212614
rect 66954 176614 67574 212058
rect 66954 176058 66986 176614
rect 67542 176058 67574 176614
rect 66954 140614 67574 176058
rect 66954 140058 66986 140614
rect 67542 140058 67574 140614
rect 66954 104614 67574 140058
rect 66954 104058 66986 104614
rect 67542 104058 67574 104614
rect 66954 68614 67574 104058
rect 66954 68058 66986 68614
rect 67542 68058 67574 68614
rect 66954 32614 67574 68058
rect 66954 32058 66986 32614
rect 67542 32058 67574 32614
rect 48954 -6662 48986 -6106
rect 49542 -6662 49574 -6106
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704282 73826 704838
rect 74382 704282 74414 704838
rect 73794 687454 74414 704282
rect 73794 686898 73826 687454
rect 74382 686898 74414 687454
rect 73794 651454 74414 686898
rect 73794 650898 73826 651454
rect 74382 650898 74414 651454
rect 73794 615454 74414 650898
rect 73794 614898 73826 615454
rect 74382 614898 74414 615454
rect 73794 579454 74414 614898
rect 73794 578898 73826 579454
rect 74382 578898 74414 579454
rect 73794 543454 74414 578898
rect 73794 542898 73826 543454
rect 74382 542898 74414 543454
rect 73794 507454 74414 542898
rect 73794 506898 73826 507454
rect 74382 506898 74414 507454
rect 73794 471454 74414 506898
rect 73794 470898 73826 471454
rect 74382 470898 74414 471454
rect 73794 435454 74414 470898
rect 73794 434898 73826 435454
rect 74382 434898 74414 435454
rect 73794 399454 74414 434898
rect 73794 398898 73826 399454
rect 74382 398898 74414 399454
rect 73794 363454 74414 398898
rect 73794 362898 73826 363454
rect 74382 362898 74414 363454
rect 73794 327454 74414 362898
rect 73794 326898 73826 327454
rect 74382 326898 74414 327454
rect 73794 291454 74414 326898
rect 73794 290898 73826 291454
rect 74382 290898 74414 291454
rect 73794 255454 74414 290898
rect 73794 254898 73826 255454
rect 74382 254898 74414 255454
rect 73794 219454 74414 254898
rect 73794 218898 73826 219454
rect 74382 218898 74414 219454
rect 73794 183454 74414 218898
rect 73794 182898 73826 183454
rect 74382 182898 74414 183454
rect 73794 147454 74414 182898
rect 73794 146898 73826 147454
rect 74382 146898 74414 147454
rect 73794 111454 74414 146898
rect 73794 110898 73826 111454
rect 74382 110898 74414 111454
rect 73794 75454 74414 110898
rect 73794 74898 73826 75454
rect 74382 74898 74414 75454
rect 73794 39454 74414 74898
rect 73794 38898 73826 39454
rect 74382 38898 74414 39454
rect 73794 3454 74414 38898
rect 73794 2898 73826 3454
rect 74382 2898 74414 3454
rect 73794 -346 74414 2898
rect 73794 -902 73826 -346
rect 74382 -902 74414 -346
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690618 77546 691174
rect 78102 690618 78134 691174
rect 77514 655174 78134 690618
rect 77514 654618 77546 655174
rect 78102 654618 78134 655174
rect 77514 619174 78134 654618
rect 77514 618618 77546 619174
rect 78102 618618 78134 619174
rect 77514 583174 78134 618618
rect 77514 582618 77546 583174
rect 78102 582618 78134 583174
rect 77514 547174 78134 582618
rect 77514 546618 77546 547174
rect 78102 546618 78134 547174
rect 77514 511174 78134 546618
rect 77514 510618 77546 511174
rect 78102 510618 78134 511174
rect 77514 475174 78134 510618
rect 77514 474618 77546 475174
rect 78102 474618 78134 475174
rect 77514 439174 78134 474618
rect 77514 438618 77546 439174
rect 78102 438618 78134 439174
rect 77514 403174 78134 438618
rect 77514 402618 77546 403174
rect 78102 402618 78134 403174
rect 77514 367174 78134 402618
rect 77514 366618 77546 367174
rect 78102 366618 78134 367174
rect 77514 331174 78134 366618
rect 77514 330618 77546 331174
rect 78102 330618 78134 331174
rect 77514 295174 78134 330618
rect 77514 294618 77546 295174
rect 78102 294618 78134 295174
rect 77514 259174 78134 294618
rect 77514 258618 77546 259174
rect 78102 258618 78134 259174
rect 77514 223174 78134 258618
rect 77514 222618 77546 223174
rect 78102 222618 78134 223174
rect 77514 187174 78134 222618
rect 77514 186618 77546 187174
rect 78102 186618 78134 187174
rect 77514 151174 78134 186618
rect 77514 150618 77546 151174
rect 78102 150618 78134 151174
rect 77514 115174 78134 150618
rect 77514 114618 77546 115174
rect 78102 114618 78134 115174
rect 77514 79174 78134 114618
rect 77514 78618 77546 79174
rect 78102 78618 78134 79174
rect 77514 43174 78134 78618
rect 77514 42618 77546 43174
rect 78102 42618 78134 43174
rect 77514 7174 78134 42618
rect 77514 6618 77546 7174
rect 78102 6618 78134 7174
rect 77514 -2266 78134 6618
rect 77514 -2822 77546 -2266
rect 78102 -2822 78134 -2266
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694338 81266 694894
rect 81822 694338 81854 694894
rect 81234 658894 81854 694338
rect 81234 658338 81266 658894
rect 81822 658338 81854 658894
rect 81234 622894 81854 658338
rect 81234 622338 81266 622894
rect 81822 622338 81854 622894
rect 81234 586894 81854 622338
rect 81234 586338 81266 586894
rect 81822 586338 81854 586894
rect 81234 550894 81854 586338
rect 81234 550338 81266 550894
rect 81822 550338 81854 550894
rect 81234 514894 81854 550338
rect 81234 514338 81266 514894
rect 81822 514338 81854 514894
rect 81234 478894 81854 514338
rect 81234 478338 81266 478894
rect 81822 478338 81854 478894
rect 81234 442894 81854 478338
rect 81234 442338 81266 442894
rect 81822 442338 81854 442894
rect 81234 406894 81854 442338
rect 81234 406338 81266 406894
rect 81822 406338 81854 406894
rect 81234 370894 81854 406338
rect 81234 370338 81266 370894
rect 81822 370338 81854 370894
rect 81234 334894 81854 370338
rect 81234 334338 81266 334894
rect 81822 334338 81854 334894
rect 81234 298894 81854 334338
rect 81234 298338 81266 298894
rect 81822 298338 81854 298894
rect 81234 262894 81854 298338
rect 81234 262338 81266 262894
rect 81822 262338 81854 262894
rect 81234 226894 81854 262338
rect 81234 226338 81266 226894
rect 81822 226338 81854 226894
rect 81234 190894 81854 226338
rect 81234 190338 81266 190894
rect 81822 190338 81854 190894
rect 81234 154894 81854 190338
rect 81234 154338 81266 154894
rect 81822 154338 81854 154894
rect 81234 118894 81854 154338
rect 81234 118338 81266 118894
rect 81822 118338 81854 118894
rect 81234 82894 81854 118338
rect 81234 82338 81266 82894
rect 81822 82338 81854 82894
rect 81234 46894 81854 82338
rect 81234 46338 81266 46894
rect 81822 46338 81854 46894
rect 81234 10894 81854 46338
rect 81234 10338 81266 10894
rect 81822 10338 81854 10894
rect 81234 -4186 81854 10338
rect 81234 -4742 81266 -4186
rect 81822 -4742 81854 -4186
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711002 102986 711558
rect 103542 711002 103574 711558
rect 99234 709638 99854 709670
rect 99234 709082 99266 709638
rect 99822 709082 99854 709638
rect 95514 707718 96134 707750
rect 95514 707162 95546 707718
rect 96102 707162 96134 707718
rect 84954 698058 84986 698614
rect 85542 698058 85574 698614
rect 84954 662614 85574 698058
rect 84954 662058 84986 662614
rect 85542 662058 85574 662614
rect 84954 626614 85574 662058
rect 84954 626058 84986 626614
rect 85542 626058 85574 626614
rect 84954 590614 85574 626058
rect 84954 590058 84986 590614
rect 85542 590058 85574 590614
rect 84954 554614 85574 590058
rect 84954 554058 84986 554614
rect 85542 554058 85574 554614
rect 84954 518614 85574 554058
rect 84954 518058 84986 518614
rect 85542 518058 85574 518614
rect 84954 482614 85574 518058
rect 84954 482058 84986 482614
rect 85542 482058 85574 482614
rect 84954 446614 85574 482058
rect 84954 446058 84986 446614
rect 85542 446058 85574 446614
rect 84954 410614 85574 446058
rect 84954 410058 84986 410614
rect 85542 410058 85574 410614
rect 84954 374614 85574 410058
rect 84954 374058 84986 374614
rect 85542 374058 85574 374614
rect 84954 338614 85574 374058
rect 84954 338058 84986 338614
rect 85542 338058 85574 338614
rect 84954 302614 85574 338058
rect 84954 302058 84986 302614
rect 85542 302058 85574 302614
rect 84954 266614 85574 302058
rect 84954 266058 84986 266614
rect 85542 266058 85574 266614
rect 84954 230614 85574 266058
rect 84954 230058 84986 230614
rect 85542 230058 85574 230614
rect 84954 194614 85574 230058
rect 84954 194058 84986 194614
rect 85542 194058 85574 194614
rect 84954 158614 85574 194058
rect 84954 158058 84986 158614
rect 85542 158058 85574 158614
rect 84954 122614 85574 158058
rect 84954 122058 84986 122614
rect 85542 122058 85574 122614
rect 84954 86614 85574 122058
rect 84954 86058 84986 86614
rect 85542 86058 85574 86614
rect 84954 50614 85574 86058
rect 84954 50058 84986 50614
rect 85542 50058 85574 50614
rect 84954 14614 85574 50058
rect 84954 14058 84986 14614
rect 85542 14058 85574 14614
rect 66954 -7622 66986 -7066
rect 67542 -7622 67574 -7066
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705242 91826 705798
rect 92382 705242 92414 705798
rect 91794 669454 92414 705242
rect 91794 668898 91826 669454
rect 92382 668898 92414 669454
rect 91794 633454 92414 668898
rect 91794 632898 91826 633454
rect 92382 632898 92414 633454
rect 91794 597454 92414 632898
rect 91794 596898 91826 597454
rect 92382 596898 92414 597454
rect 91794 561454 92414 596898
rect 91794 560898 91826 561454
rect 92382 560898 92414 561454
rect 91794 525454 92414 560898
rect 91794 524898 91826 525454
rect 92382 524898 92414 525454
rect 91794 489454 92414 524898
rect 91794 488898 91826 489454
rect 92382 488898 92414 489454
rect 91794 453454 92414 488898
rect 91794 452898 91826 453454
rect 92382 452898 92414 453454
rect 91794 417454 92414 452898
rect 91794 416898 91826 417454
rect 92382 416898 92414 417454
rect 91794 381454 92414 416898
rect 91794 380898 91826 381454
rect 92382 380898 92414 381454
rect 91794 345454 92414 380898
rect 91794 344898 91826 345454
rect 92382 344898 92414 345454
rect 91794 309454 92414 344898
rect 91794 308898 91826 309454
rect 92382 308898 92414 309454
rect 91794 273454 92414 308898
rect 91794 272898 91826 273454
rect 92382 272898 92414 273454
rect 91794 237454 92414 272898
rect 91794 236898 91826 237454
rect 92382 236898 92414 237454
rect 91794 201454 92414 236898
rect 91794 200898 91826 201454
rect 92382 200898 92414 201454
rect 91794 165454 92414 200898
rect 91794 164898 91826 165454
rect 92382 164898 92414 165454
rect 91794 129454 92414 164898
rect 91794 128898 91826 129454
rect 92382 128898 92414 129454
rect 91794 93454 92414 128898
rect 91794 92898 91826 93454
rect 92382 92898 92414 93454
rect 91794 57454 92414 92898
rect 91794 56898 91826 57454
rect 92382 56898 92414 57454
rect 91794 21454 92414 56898
rect 91794 20898 91826 21454
rect 92382 20898 92414 21454
rect 91794 -1306 92414 20898
rect 91794 -1862 91826 -1306
rect 92382 -1862 92414 -1306
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672618 95546 673174
rect 96102 672618 96134 673174
rect 95514 637174 96134 672618
rect 95514 636618 95546 637174
rect 96102 636618 96134 637174
rect 95514 601174 96134 636618
rect 95514 600618 95546 601174
rect 96102 600618 96134 601174
rect 95514 565174 96134 600618
rect 95514 564618 95546 565174
rect 96102 564618 96134 565174
rect 95514 529174 96134 564618
rect 95514 528618 95546 529174
rect 96102 528618 96134 529174
rect 95514 493174 96134 528618
rect 95514 492618 95546 493174
rect 96102 492618 96134 493174
rect 95514 457174 96134 492618
rect 95514 456618 95546 457174
rect 96102 456618 96134 457174
rect 95514 421174 96134 456618
rect 95514 420618 95546 421174
rect 96102 420618 96134 421174
rect 95514 385174 96134 420618
rect 95514 384618 95546 385174
rect 96102 384618 96134 385174
rect 95514 349174 96134 384618
rect 95514 348618 95546 349174
rect 96102 348618 96134 349174
rect 95514 313174 96134 348618
rect 95514 312618 95546 313174
rect 96102 312618 96134 313174
rect 95514 277174 96134 312618
rect 95514 276618 95546 277174
rect 96102 276618 96134 277174
rect 95514 241174 96134 276618
rect 95514 240618 95546 241174
rect 96102 240618 96134 241174
rect 95514 205174 96134 240618
rect 95514 204618 95546 205174
rect 96102 204618 96134 205174
rect 95514 169174 96134 204618
rect 95514 168618 95546 169174
rect 96102 168618 96134 169174
rect 95514 133174 96134 168618
rect 95514 132618 95546 133174
rect 96102 132618 96134 133174
rect 95514 97174 96134 132618
rect 95514 96618 95546 97174
rect 96102 96618 96134 97174
rect 95514 61174 96134 96618
rect 95514 60618 95546 61174
rect 96102 60618 96134 61174
rect 95514 25174 96134 60618
rect 95514 24618 95546 25174
rect 96102 24618 96134 25174
rect 95514 -3226 96134 24618
rect 95514 -3782 95546 -3226
rect 96102 -3782 96134 -3226
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676338 99266 676894
rect 99822 676338 99854 676894
rect 99234 640894 99854 676338
rect 99234 640338 99266 640894
rect 99822 640338 99854 640894
rect 99234 604894 99854 640338
rect 99234 604338 99266 604894
rect 99822 604338 99854 604894
rect 99234 568894 99854 604338
rect 99234 568338 99266 568894
rect 99822 568338 99854 568894
rect 99234 532894 99854 568338
rect 99234 532338 99266 532894
rect 99822 532338 99854 532894
rect 99234 496894 99854 532338
rect 99234 496338 99266 496894
rect 99822 496338 99854 496894
rect 99234 460894 99854 496338
rect 99234 460338 99266 460894
rect 99822 460338 99854 460894
rect 99234 424894 99854 460338
rect 99234 424338 99266 424894
rect 99822 424338 99854 424894
rect 99234 388894 99854 424338
rect 99234 388338 99266 388894
rect 99822 388338 99854 388894
rect 99234 352894 99854 388338
rect 99234 352338 99266 352894
rect 99822 352338 99854 352894
rect 99234 316894 99854 352338
rect 99234 316338 99266 316894
rect 99822 316338 99854 316894
rect 99234 280894 99854 316338
rect 99234 280338 99266 280894
rect 99822 280338 99854 280894
rect 99234 244894 99854 280338
rect 99234 244338 99266 244894
rect 99822 244338 99854 244894
rect 99234 208894 99854 244338
rect 99234 208338 99266 208894
rect 99822 208338 99854 208894
rect 99234 172894 99854 208338
rect 99234 172338 99266 172894
rect 99822 172338 99854 172894
rect 99234 136894 99854 172338
rect 99234 136338 99266 136894
rect 99822 136338 99854 136894
rect 99234 100894 99854 136338
rect 99234 100338 99266 100894
rect 99822 100338 99854 100894
rect 99234 64894 99854 100338
rect 99234 64338 99266 64894
rect 99822 64338 99854 64894
rect 99234 28894 99854 64338
rect 99234 28338 99266 28894
rect 99822 28338 99854 28894
rect 99234 -5146 99854 28338
rect 99234 -5702 99266 -5146
rect 99822 -5702 99854 -5146
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710042 120986 710598
rect 121542 710042 121574 710598
rect 117234 708678 117854 709670
rect 117234 708122 117266 708678
rect 117822 708122 117854 708678
rect 113514 706758 114134 707750
rect 113514 706202 113546 706758
rect 114102 706202 114134 706758
rect 102954 680058 102986 680614
rect 103542 680058 103574 680614
rect 102954 644614 103574 680058
rect 102954 644058 102986 644614
rect 103542 644058 103574 644614
rect 102954 608614 103574 644058
rect 102954 608058 102986 608614
rect 103542 608058 103574 608614
rect 102954 572614 103574 608058
rect 102954 572058 102986 572614
rect 103542 572058 103574 572614
rect 102954 536614 103574 572058
rect 102954 536058 102986 536614
rect 103542 536058 103574 536614
rect 102954 500614 103574 536058
rect 102954 500058 102986 500614
rect 103542 500058 103574 500614
rect 102954 464614 103574 500058
rect 102954 464058 102986 464614
rect 103542 464058 103574 464614
rect 102954 428614 103574 464058
rect 102954 428058 102986 428614
rect 103542 428058 103574 428614
rect 102954 392614 103574 428058
rect 102954 392058 102986 392614
rect 103542 392058 103574 392614
rect 102954 356614 103574 392058
rect 102954 356058 102986 356614
rect 103542 356058 103574 356614
rect 102954 320614 103574 356058
rect 102954 320058 102986 320614
rect 103542 320058 103574 320614
rect 102954 284614 103574 320058
rect 102954 284058 102986 284614
rect 103542 284058 103574 284614
rect 102954 248614 103574 284058
rect 102954 248058 102986 248614
rect 103542 248058 103574 248614
rect 102954 212614 103574 248058
rect 102954 212058 102986 212614
rect 103542 212058 103574 212614
rect 102954 176614 103574 212058
rect 102954 176058 102986 176614
rect 103542 176058 103574 176614
rect 102954 140614 103574 176058
rect 102954 140058 102986 140614
rect 103542 140058 103574 140614
rect 102954 104614 103574 140058
rect 102954 104058 102986 104614
rect 103542 104058 103574 104614
rect 102954 68614 103574 104058
rect 102954 68058 102986 68614
rect 103542 68058 103574 68614
rect 102954 32614 103574 68058
rect 102954 32058 102986 32614
rect 103542 32058 103574 32614
rect 84954 -6662 84986 -6106
rect 85542 -6662 85574 -6106
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704282 109826 704838
rect 110382 704282 110414 704838
rect 109794 687454 110414 704282
rect 109794 686898 109826 687454
rect 110382 686898 110414 687454
rect 109794 651454 110414 686898
rect 109794 650898 109826 651454
rect 110382 650898 110414 651454
rect 109794 615454 110414 650898
rect 109794 614898 109826 615454
rect 110382 614898 110414 615454
rect 109794 579454 110414 614898
rect 109794 578898 109826 579454
rect 110382 578898 110414 579454
rect 109794 543454 110414 578898
rect 109794 542898 109826 543454
rect 110382 542898 110414 543454
rect 109794 507454 110414 542898
rect 109794 506898 109826 507454
rect 110382 506898 110414 507454
rect 109794 471454 110414 506898
rect 109794 470898 109826 471454
rect 110382 470898 110414 471454
rect 109794 435454 110414 470898
rect 109794 434898 109826 435454
rect 110382 434898 110414 435454
rect 109794 399454 110414 434898
rect 109794 398898 109826 399454
rect 110382 398898 110414 399454
rect 109794 363454 110414 398898
rect 109794 362898 109826 363454
rect 110382 362898 110414 363454
rect 109794 327454 110414 362898
rect 109794 326898 109826 327454
rect 110382 326898 110414 327454
rect 109794 291454 110414 326898
rect 109794 290898 109826 291454
rect 110382 290898 110414 291454
rect 109794 255454 110414 290898
rect 109794 254898 109826 255454
rect 110382 254898 110414 255454
rect 109794 219454 110414 254898
rect 109794 218898 109826 219454
rect 110382 218898 110414 219454
rect 109794 183454 110414 218898
rect 109794 182898 109826 183454
rect 110382 182898 110414 183454
rect 109794 147454 110414 182898
rect 109794 146898 109826 147454
rect 110382 146898 110414 147454
rect 109794 111454 110414 146898
rect 109794 110898 109826 111454
rect 110382 110898 110414 111454
rect 109794 75454 110414 110898
rect 109794 74898 109826 75454
rect 110382 74898 110414 75454
rect 109794 39454 110414 74898
rect 109794 38898 109826 39454
rect 110382 38898 110414 39454
rect 109794 3454 110414 38898
rect 109794 2898 109826 3454
rect 110382 2898 110414 3454
rect 109794 -346 110414 2898
rect 109794 -902 109826 -346
rect 110382 -902 110414 -346
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690618 113546 691174
rect 114102 690618 114134 691174
rect 113514 655174 114134 690618
rect 113514 654618 113546 655174
rect 114102 654618 114134 655174
rect 113514 619174 114134 654618
rect 113514 618618 113546 619174
rect 114102 618618 114134 619174
rect 113514 583174 114134 618618
rect 113514 582618 113546 583174
rect 114102 582618 114134 583174
rect 113514 547174 114134 582618
rect 113514 546618 113546 547174
rect 114102 546618 114134 547174
rect 113514 511174 114134 546618
rect 113514 510618 113546 511174
rect 114102 510618 114134 511174
rect 113514 475174 114134 510618
rect 113514 474618 113546 475174
rect 114102 474618 114134 475174
rect 113514 439174 114134 474618
rect 113514 438618 113546 439174
rect 114102 438618 114134 439174
rect 113514 403174 114134 438618
rect 113514 402618 113546 403174
rect 114102 402618 114134 403174
rect 113514 367174 114134 402618
rect 113514 366618 113546 367174
rect 114102 366618 114134 367174
rect 113514 331174 114134 366618
rect 113514 330618 113546 331174
rect 114102 330618 114134 331174
rect 113514 295174 114134 330618
rect 113514 294618 113546 295174
rect 114102 294618 114134 295174
rect 113514 259174 114134 294618
rect 113514 258618 113546 259174
rect 114102 258618 114134 259174
rect 113514 223174 114134 258618
rect 113514 222618 113546 223174
rect 114102 222618 114134 223174
rect 113514 187174 114134 222618
rect 113514 186618 113546 187174
rect 114102 186618 114134 187174
rect 113514 151174 114134 186618
rect 113514 150618 113546 151174
rect 114102 150618 114134 151174
rect 113514 115174 114134 150618
rect 113514 114618 113546 115174
rect 114102 114618 114134 115174
rect 113514 79174 114134 114618
rect 113514 78618 113546 79174
rect 114102 78618 114134 79174
rect 113514 43174 114134 78618
rect 113514 42618 113546 43174
rect 114102 42618 114134 43174
rect 113514 7174 114134 42618
rect 113514 6618 113546 7174
rect 114102 6618 114134 7174
rect 113514 -2266 114134 6618
rect 113514 -2822 113546 -2266
rect 114102 -2822 114134 -2266
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694338 117266 694894
rect 117822 694338 117854 694894
rect 117234 658894 117854 694338
rect 117234 658338 117266 658894
rect 117822 658338 117854 658894
rect 117234 622894 117854 658338
rect 117234 622338 117266 622894
rect 117822 622338 117854 622894
rect 117234 586894 117854 622338
rect 117234 586338 117266 586894
rect 117822 586338 117854 586894
rect 117234 550894 117854 586338
rect 117234 550338 117266 550894
rect 117822 550338 117854 550894
rect 117234 514894 117854 550338
rect 117234 514338 117266 514894
rect 117822 514338 117854 514894
rect 117234 478894 117854 514338
rect 117234 478338 117266 478894
rect 117822 478338 117854 478894
rect 117234 442894 117854 478338
rect 117234 442338 117266 442894
rect 117822 442338 117854 442894
rect 117234 406894 117854 442338
rect 117234 406338 117266 406894
rect 117822 406338 117854 406894
rect 117234 370894 117854 406338
rect 117234 370338 117266 370894
rect 117822 370338 117854 370894
rect 117234 334894 117854 370338
rect 117234 334338 117266 334894
rect 117822 334338 117854 334894
rect 117234 298894 117854 334338
rect 117234 298338 117266 298894
rect 117822 298338 117854 298894
rect 117234 262894 117854 298338
rect 117234 262338 117266 262894
rect 117822 262338 117854 262894
rect 117234 226894 117854 262338
rect 117234 226338 117266 226894
rect 117822 226338 117854 226894
rect 117234 190894 117854 226338
rect 117234 190338 117266 190894
rect 117822 190338 117854 190894
rect 117234 154894 117854 190338
rect 117234 154338 117266 154894
rect 117822 154338 117854 154894
rect 117234 118894 117854 154338
rect 117234 118338 117266 118894
rect 117822 118338 117854 118894
rect 117234 82894 117854 118338
rect 117234 82338 117266 82894
rect 117822 82338 117854 82894
rect 117234 46894 117854 82338
rect 117234 46338 117266 46894
rect 117822 46338 117854 46894
rect 117234 10894 117854 46338
rect 117234 10338 117266 10894
rect 117822 10338 117854 10894
rect 117234 -4186 117854 10338
rect 117234 -4742 117266 -4186
rect 117822 -4742 117854 -4186
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711002 138986 711558
rect 139542 711002 139574 711558
rect 135234 709638 135854 709670
rect 135234 709082 135266 709638
rect 135822 709082 135854 709638
rect 131514 707718 132134 707750
rect 131514 707162 131546 707718
rect 132102 707162 132134 707718
rect 120954 698058 120986 698614
rect 121542 698058 121574 698614
rect 120954 662614 121574 698058
rect 120954 662058 120986 662614
rect 121542 662058 121574 662614
rect 120954 626614 121574 662058
rect 120954 626058 120986 626614
rect 121542 626058 121574 626614
rect 120954 590614 121574 626058
rect 120954 590058 120986 590614
rect 121542 590058 121574 590614
rect 120954 554614 121574 590058
rect 120954 554058 120986 554614
rect 121542 554058 121574 554614
rect 120954 518614 121574 554058
rect 120954 518058 120986 518614
rect 121542 518058 121574 518614
rect 120954 482614 121574 518058
rect 120954 482058 120986 482614
rect 121542 482058 121574 482614
rect 120954 446614 121574 482058
rect 120954 446058 120986 446614
rect 121542 446058 121574 446614
rect 120954 410614 121574 446058
rect 120954 410058 120986 410614
rect 121542 410058 121574 410614
rect 120954 374614 121574 410058
rect 120954 374058 120986 374614
rect 121542 374058 121574 374614
rect 120954 338614 121574 374058
rect 120954 338058 120986 338614
rect 121542 338058 121574 338614
rect 120954 302614 121574 338058
rect 120954 302058 120986 302614
rect 121542 302058 121574 302614
rect 120954 266614 121574 302058
rect 120954 266058 120986 266614
rect 121542 266058 121574 266614
rect 120954 230614 121574 266058
rect 120954 230058 120986 230614
rect 121542 230058 121574 230614
rect 120954 194614 121574 230058
rect 120954 194058 120986 194614
rect 121542 194058 121574 194614
rect 120954 158614 121574 194058
rect 120954 158058 120986 158614
rect 121542 158058 121574 158614
rect 120954 122614 121574 158058
rect 120954 122058 120986 122614
rect 121542 122058 121574 122614
rect 120954 86614 121574 122058
rect 120954 86058 120986 86614
rect 121542 86058 121574 86614
rect 120954 50614 121574 86058
rect 120954 50058 120986 50614
rect 121542 50058 121574 50614
rect 120954 14614 121574 50058
rect 120954 14058 120986 14614
rect 121542 14058 121574 14614
rect 102954 -7622 102986 -7066
rect 103542 -7622 103574 -7066
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705242 127826 705798
rect 128382 705242 128414 705798
rect 127794 669454 128414 705242
rect 127794 668898 127826 669454
rect 128382 668898 128414 669454
rect 127794 633454 128414 668898
rect 127794 632898 127826 633454
rect 128382 632898 128414 633454
rect 127794 597454 128414 632898
rect 127794 596898 127826 597454
rect 128382 596898 128414 597454
rect 127794 561454 128414 596898
rect 127794 560898 127826 561454
rect 128382 560898 128414 561454
rect 127794 525454 128414 560898
rect 127794 524898 127826 525454
rect 128382 524898 128414 525454
rect 127794 489454 128414 524898
rect 127794 488898 127826 489454
rect 128382 488898 128414 489454
rect 127794 453454 128414 488898
rect 127794 452898 127826 453454
rect 128382 452898 128414 453454
rect 127794 417454 128414 452898
rect 127794 416898 127826 417454
rect 128382 416898 128414 417454
rect 127794 381454 128414 416898
rect 127794 380898 127826 381454
rect 128382 380898 128414 381454
rect 127794 345454 128414 380898
rect 127794 344898 127826 345454
rect 128382 344898 128414 345454
rect 127794 309454 128414 344898
rect 127794 308898 127826 309454
rect 128382 308898 128414 309454
rect 127794 273454 128414 308898
rect 127794 272898 127826 273454
rect 128382 272898 128414 273454
rect 127794 237454 128414 272898
rect 127794 236898 127826 237454
rect 128382 236898 128414 237454
rect 127794 201454 128414 236898
rect 127794 200898 127826 201454
rect 128382 200898 128414 201454
rect 127794 165454 128414 200898
rect 127794 164898 127826 165454
rect 128382 164898 128414 165454
rect 127794 129454 128414 164898
rect 127794 128898 127826 129454
rect 128382 128898 128414 129454
rect 127794 93454 128414 128898
rect 127794 92898 127826 93454
rect 128382 92898 128414 93454
rect 127794 57454 128414 92898
rect 127794 56898 127826 57454
rect 128382 56898 128414 57454
rect 127794 21454 128414 56898
rect 127794 20898 127826 21454
rect 128382 20898 128414 21454
rect 127794 -1306 128414 20898
rect 127794 -1862 127826 -1306
rect 128382 -1862 128414 -1306
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672618 131546 673174
rect 132102 672618 132134 673174
rect 131514 637174 132134 672618
rect 131514 636618 131546 637174
rect 132102 636618 132134 637174
rect 131514 601174 132134 636618
rect 131514 600618 131546 601174
rect 132102 600618 132134 601174
rect 131514 565174 132134 600618
rect 131514 564618 131546 565174
rect 132102 564618 132134 565174
rect 131514 529174 132134 564618
rect 131514 528618 131546 529174
rect 132102 528618 132134 529174
rect 131514 493174 132134 528618
rect 131514 492618 131546 493174
rect 132102 492618 132134 493174
rect 131514 457174 132134 492618
rect 131514 456618 131546 457174
rect 132102 456618 132134 457174
rect 131514 421174 132134 456618
rect 131514 420618 131546 421174
rect 132102 420618 132134 421174
rect 131514 385174 132134 420618
rect 131514 384618 131546 385174
rect 132102 384618 132134 385174
rect 131514 349174 132134 384618
rect 131514 348618 131546 349174
rect 132102 348618 132134 349174
rect 131514 313174 132134 348618
rect 131514 312618 131546 313174
rect 132102 312618 132134 313174
rect 131514 277174 132134 312618
rect 131514 276618 131546 277174
rect 132102 276618 132134 277174
rect 131514 241174 132134 276618
rect 131514 240618 131546 241174
rect 132102 240618 132134 241174
rect 131514 205174 132134 240618
rect 131514 204618 131546 205174
rect 132102 204618 132134 205174
rect 131514 169174 132134 204618
rect 131514 168618 131546 169174
rect 132102 168618 132134 169174
rect 131514 133174 132134 168618
rect 131514 132618 131546 133174
rect 132102 132618 132134 133174
rect 131514 97174 132134 132618
rect 131514 96618 131546 97174
rect 132102 96618 132134 97174
rect 131514 61174 132134 96618
rect 131514 60618 131546 61174
rect 132102 60618 132134 61174
rect 131514 25174 132134 60618
rect 131514 24618 131546 25174
rect 132102 24618 132134 25174
rect 131514 -3226 132134 24618
rect 131514 -3782 131546 -3226
rect 132102 -3782 132134 -3226
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676338 135266 676894
rect 135822 676338 135854 676894
rect 135234 640894 135854 676338
rect 135234 640338 135266 640894
rect 135822 640338 135854 640894
rect 135234 604894 135854 640338
rect 135234 604338 135266 604894
rect 135822 604338 135854 604894
rect 135234 568894 135854 604338
rect 135234 568338 135266 568894
rect 135822 568338 135854 568894
rect 135234 532894 135854 568338
rect 135234 532338 135266 532894
rect 135822 532338 135854 532894
rect 135234 496894 135854 532338
rect 135234 496338 135266 496894
rect 135822 496338 135854 496894
rect 135234 460894 135854 496338
rect 135234 460338 135266 460894
rect 135822 460338 135854 460894
rect 135234 424894 135854 460338
rect 135234 424338 135266 424894
rect 135822 424338 135854 424894
rect 135234 388894 135854 424338
rect 135234 388338 135266 388894
rect 135822 388338 135854 388894
rect 135234 352894 135854 388338
rect 135234 352338 135266 352894
rect 135822 352338 135854 352894
rect 135234 316894 135854 352338
rect 135234 316338 135266 316894
rect 135822 316338 135854 316894
rect 135234 280894 135854 316338
rect 135234 280338 135266 280894
rect 135822 280338 135854 280894
rect 135234 244894 135854 280338
rect 135234 244338 135266 244894
rect 135822 244338 135854 244894
rect 135234 208894 135854 244338
rect 135234 208338 135266 208894
rect 135822 208338 135854 208894
rect 135234 172894 135854 208338
rect 135234 172338 135266 172894
rect 135822 172338 135854 172894
rect 135234 136894 135854 172338
rect 135234 136338 135266 136894
rect 135822 136338 135854 136894
rect 135234 100894 135854 136338
rect 135234 100338 135266 100894
rect 135822 100338 135854 100894
rect 135234 64894 135854 100338
rect 135234 64338 135266 64894
rect 135822 64338 135854 64894
rect 135234 28894 135854 64338
rect 135234 28338 135266 28894
rect 135822 28338 135854 28894
rect 135234 -5146 135854 28338
rect 135234 -5702 135266 -5146
rect 135822 -5702 135854 -5146
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710042 156986 710598
rect 157542 710042 157574 710598
rect 153234 708678 153854 709670
rect 153234 708122 153266 708678
rect 153822 708122 153854 708678
rect 149514 706758 150134 707750
rect 149514 706202 149546 706758
rect 150102 706202 150134 706758
rect 138954 680058 138986 680614
rect 139542 680058 139574 680614
rect 138954 644614 139574 680058
rect 138954 644058 138986 644614
rect 139542 644058 139574 644614
rect 138954 608614 139574 644058
rect 138954 608058 138986 608614
rect 139542 608058 139574 608614
rect 138954 572614 139574 608058
rect 138954 572058 138986 572614
rect 139542 572058 139574 572614
rect 138954 536614 139574 572058
rect 138954 536058 138986 536614
rect 139542 536058 139574 536614
rect 138954 500614 139574 536058
rect 138954 500058 138986 500614
rect 139542 500058 139574 500614
rect 138954 464614 139574 500058
rect 138954 464058 138986 464614
rect 139542 464058 139574 464614
rect 138954 428614 139574 464058
rect 138954 428058 138986 428614
rect 139542 428058 139574 428614
rect 138954 392614 139574 428058
rect 138954 392058 138986 392614
rect 139542 392058 139574 392614
rect 138954 356614 139574 392058
rect 138954 356058 138986 356614
rect 139542 356058 139574 356614
rect 138954 320614 139574 356058
rect 138954 320058 138986 320614
rect 139542 320058 139574 320614
rect 138954 284614 139574 320058
rect 138954 284058 138986 284614
rect 139542 284058 139574 284614
rect 138954 248614 139574 284058
rect 138954 248058 138986 248614
rect 139542 248058 139574 248614
rect 138954 212614 139574 248058
rect 138954 212058 138986 212614
rect 139542 212058 139574 212614
rect 138954 176614 139574 212058
rect 138954 176058 138986 176614
rect 139542 176058 139574 176614
rect 138954 140614 139574 176058
rect 138954 140058 138986 140614
rect 139542 140058 139574 140614
rect 138954 104614 139574 140058
rect 138954 104058 138986 104614
rect 139542 104058 139574 104614
rect 138954 68614 139574 104058
rect 138954 68058 138986 68614
rect 139542 68058 139574 68614
rect 138954 32614 139574 68058
rect 138954 32058 138986 32614
rect 139542 32058 139574 32614
rect 120954 -6662 120986 -6106
rect 121542 -6662 121574 -6106
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704282 145826 704838
rect 146382 704282 146414 704838
rect 145794 687454 146414 704282
rect 145794 686898 145826 687454
rect 146382 686898 146414 687454
rect 145794 651454 146414 686898
rect 145794 650898 145826 651454
rect 146382 650898 146414 651454
rect 145794 615454 146414 650898
rect 145794 614898 145826 615454
rect 146382 614898 146414 615454
rect 145794 579454 146414 614898
rect 145794 578898 145826 579454
rect 146382 578898 146414 579454
rect 145794 543454 146414 578898
rect 145794 542898 145826 543454
rect 146382 542898 146414 543454
rect 145794 507454 146414 542898
rect 145794 506898 145826 507454
rect 146382 506898 146414 507454
rect 145794 471454 146414 506898
rect 145794 470898 145826 471454
rect 146382 470898 146414 471454
rect 145794 435454 146414 470898
rect 145794 434898 145826 435454
rect 146382 434898 146414 435454
rect 145794 399454 146414 434898
rect 145794 398898 145826 399454
rect 146382 398898 146414 399454
rect 145794 363454 146414 398898
rect 145794 362898 145826 363454
rect 146382 362898 146414 363454
rect 145794 327454 146414 362898
rect 145794 326898 145826 327454
rect 146382 326898 146414 327454
rect 145794 291454 146414 326898
rect 145794 290898 145826 291454
rect 146382 290898 146414 291454
rect 145794 255454 146414 290898
rect 145794 254898 145826 255454
rect 146382 254898 146414 255454
rect 145794 219454 146414 254898
rect 145794 218898 145826 219454
rect 146382 218898 146414 219454
rect 145794 183454 146414 218898
rect 145794 182898 145826 183454
rect 146382 182898 146414 183454
rect 145794 147454 146414 182898
rect 145794 146898 145826 147454
rect 146382 146898 146414 147454
rect 145794 111454 146414 146898
rect 145794 110898 145826 111454
rect 146382 110898 146414 111454
rect 145794 75454 146414 110898
rect 145794 74898 145826 75454
rect 146382 74898 146414 75454
rect 145794 39454 146414 74898
rect 145794 38898 145826 39454
rect 146382 38898 146414 39454
rect 145794 3454 146414 38898
rect 145794 2898 145826 3454
rect 146382 2898 146414 3454
rect 145794 -346 146414 2898
rect 145794 -902 145826 -346
rect 146382 -902 146414 -346
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690618 149546 691174
rect 150102 690618 150134 691174
rect 149514 655174 150134 690618
rect 149514 654618 149546 655174
rect 150102 654618 150134 655174
rect 149514 619174 150134 654618
rect 149514 618618 149546 619174
rect 150102 618618 150134 619174
rect 149514 583174 150134 618618
rect 149514 582618 149546 583174
rect 150102 582618 150134 583174
rect 149514 547174 150134 582618
rect 149514 546618 149546 547174
rect 150102 546618 150134 547174
rect 149514 511174 150134 546618
rect 149514 510618 149546 511174
rect 150102 510618 150134 511174
rect 149514 475174 150134 510618
rect 149514 474618 149546 475174
rect 150102 474618 150134 475174
rect 149514 439174 150134 474618
rect 149514 438618 149546 439174
rect 150102 438618 150134 439174
rect 149514 403174 150134 438618
rect 149514 402618 149546 403174
rect 150102 402618 150134 403174
rect 149514 367174 150134 402618
rect 149514 366618 149546 367174
rect 150102 366618 150134 367174
rect 149514 331174 150134 366618
rect 149514 330618 149546 331174
rect 150102 330618 150134 331174
rect 149514 295174 150134 330618
rect 149514 294618 149546 295174
rect 150102 294618 150134 295174
rect 149514 259174 150134 294618
rect 149514 258618 149546 259174
rect 150102 258618 150134 259174
rect 149514 223174 150134 258618
rect 149514 222618 149546 223174
rect 150102 222618 150134 223174
rect 149514 187174 150134 222618
rect 149514 186618 149546 187174
rect 150102 186618 150134 187174
rect 149514 151174 150134 186618
rect 149514 150618 149546 151174
rect 150102 150618 150134 151174
rect 149514 115174 150134 150618
rect 149514 114618 149546 115174
rect 150102 114618 150134 115174
rect 149514 79174 150134 114618
rect 149514 78618 149546 79174
rect 150102 78618 150134 79174
rect 149514 43174 150134 78618
rect 149514 42618 149546 43174
rect 150102 42618 150134 43174
rect 149514 7174 150134 42618
rect 149514 6618 149546 7174
rect 150102 6618 150134 7174
rect 149514 -2266 150134 6618
rect 149514 -2822 149546 -2266
rect 150102 -2822 150134 -2266
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694338 153266 694894
rect 153822 694338 153854 694894
rect 153234 658894 153854 694338
rect 153234 658338 153266 658894
rect 153822 658338 153854 658894
rect 153234 622894 153854 658338
rect 153234 622338 153266 622894
rect 153822 622338 153854 622894
rect 153234 586894 153854 622338
rect 153234 586338 153266 586894
rect 153822 586338 153854 586894
rect 153234 550894 153854 586338
rect 153234 550338 153266 550894
rect 153822 550338 153854 550894
rect 153234 514894 153854 550338
rect 153234 514338 153266 514894
rect 153822 514338 153854 514894
rect 153234 478894 153854 514338
rect 153234 478338 153266 478894
rect 153822 478338 153854 478894
rect 153234 442894 153854 478338
rect 153234 442338 153266 442894
rect 153822 442338 153854 442894
rect 153234 406894 153854 442338
rect 153234 406338 153266 406894
rect 153822 406338 153854 406894
rect 153234 370894 153854 406338
rect 153234 370338 153266 370894
rect 153822 370338 153854 370894
rect 153234 334894 153854 370338
rect 153234 334338 153266 334894
rect 153822 334338 153854 334894
rect 153234 298894 153854 334338
rect 153234 298338 153266 298894
rect 153822 298338 153854 298894
rect 153234 262894 153854 298338
rect 153234 262338 153266 262894
rect 153822 262338 153854 262894
rect 153234 226894 153854 262338
rect 153234 226338 153266 226894
rect 153822 226338 153854 226894
rect 153234 190894 153854 226338
rect 153234 190338 153266 190894
rect 153822 190338 153854 190894
rect 153234 154894 153854 190338
rect 153234 154338 153266 154894
rect 153822 154338 153854 154894
rect 153234 118894 153854 154338
rect 153234 118338 153266 118894
rect 153822 118338 153854 118894
rect 153234 82894 153854 118338
rect 153234 82338 153266 82894
rect 153822 82338 153854 82894
rect 153234 46894 153854 82338
rect 153234 46338 153266 46894
rect 153822 46338 153854 46894
rect 153234 10894 153854 46338
rect 153234 10338 153266 10894
rect 153822 10338 153854 10894
rect 153234 -4186 153854 10338
rect 153234 -4742 153266 -4186
rect 153822 -4742 153854 -4186
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711002 174986 711558
rect 175542 711002 175574 711558
rect 171234 709638 171854 709670
rect 171234 709082 171266 709638
rect 171822 709082 171854 709638
rect 167514 707718 168134 707750
rect 167514 707162 167546 707718
rect 168102 707162 168134 707718
rect 156954 698058 156986 698614
rect 157542 698058 157574 698614
rect 156954 662614 157574 698058
rect 156954 662058 156986 662614
rect 157542 662058 157574 662614
rect 156954 626614 157574 662058
rect 156954 626058 156986 626614
rect 157542 626058 157574 626614
rect 156954 590614 157574 626058
rect 156954 590058 156986 590614
rect 157542 590058 157574 590614
rect 156954 554614 157574 590058
rect 156954 554058 156986 554614
rect 157542 554058 157574 554614
rect 156954 518614 157574 554058
rect 156954 518058 156986 518614
rect 157542 518058 157574 518614
rect 156954 482614 157574 518058
rect 156954 482058 156986 482614
rect 157542 482058 157574 482614
rect 156954 446614 157574 482058
rect 156954 446058 156986 446614
rect 157542 446058 157574 446614
rect 156954 410614 157574 446058
rect 156954 410058 156986 410614
rect 157542 410058 157574 410614
rect 156954 374614 157574 410058
rect 156954 374058 156986 374614
rect 157542 374058 157574 374614
rect 156954 338614 157574 374058
rect 156954 338058 156986 338614
rect 157542 338058 157574 338614
rect 156954 302614 157574 338058
rect 156954 302058 156986 302614
rect 157542 302058 157574 302614
rect 156954 266614 157574 302058
rect 156954 266058 156986 266614
rect 157542 266058 157574 266614
rect 156954 230614 157574 266058
rect 156954 230058 156986 230614
rect 157542 230058 157574 230614
rect 156954 194614 157574 230058
rect 156954 194058 156986 194614
rect 157542 194058 157574 194614
rect 156954 158614 157574 194058
rect 156954 158058 156986 158614
rect 157542 158058 157574 158614
rect 156954 122614 157574 158058
rect 156954 122058 156986 122614
rect 157542 122058 157574 122614
rect 156954 86614 157574 122058
rect 156954 86058 156986 86614
rect 157542 86058 157574 86614
rect 156954 50614 157574 86058
rect 156954 50058 156986 50614
rect 157542 50058 157574 50614
rect 156954 14614 157574 50058
rect 156954 14058 156986 14614
rect 157542 14058 157574 14614
rect 138954 -7622 138986 -7066
rect 139542 -7622 139574 -7066
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705242 163826 705798
rect 164382 705242 164414 705798
rect 163794 669454 164414 705242
rect 163794 668898 163826 669454
rect 164382 668898 164414 669454
rect 163794 633454 164414 668898
rect 163794 632898 163826 633454
rect 164382 632898 164414 633454
rect 163794 597454 164414 632898
rect 163794 596898 163826 597454
rect 164382 596898 164414 597454
rect 163794 561454 164414 596898
rect 163794 560898 163826 561454
rect 164382 560898 164414 561454
rect 163794 525454 164414 560898
rect 163794 524898 163826 525454
rect 164382 524898 164414 525454
rect 163794 489454 164414 524898
rect 163794 488898 163826 489454
rect 164382 488898 164414 489454
rect 163794 453454 164414 488898
rect 163794 452898 163826 453454
rect 164382 452898 164414 453454
rect 163794 417454 164414 452898
rect 163794 416898 163826 417454
rect 164382 416898 164414 417454
rect 163794 381454 164414 416898
rect 163794 380898 163826 381454
rect 164382 380898 164414 381454
rect 163794 345454 164414 380898
rect 163794 344898 163826 345454
rect 164382 344898 164414 345454
rect 163794 309454 164414 344898
rect 163794 308898 163826 309454
rect 164382 308898 164414 309454
rect 163794 273454 164414 308898
rect 163794 272898 163826 273454
rect 164382 272898 164414 273454
rect 163794 237454 164414 272898
rect 163794 236898 163826 237454
rect 164382 236898 164414 237454
rect 163794 201454 164414 236898
rect 163794 200898 163826 201454
rect 164382 200898 164414 201454
rect 163794 165454 164414 200898
rect 163794 164898 163826 165454
rect 164382 164898 164414 165454
rect 163794 129454 164414 164898
rect 163794 128898 163826 129454
rect 164382 128898 164414 129454
rect 163794 93454 164414 128898
rect 163794 92898 163826 93454
rect 164382 92898 164414 93454
rect 163794 57454 164414 92898
rect 163794 56898 163826 57454
rect 164382 56898 164414 57454
rect 163794 21454 164414 56898
rect 163794 20898 163826 21454
rect 164382 20898 164414 21454
rect 163794 -1306 164414 20898
rect 163794 -1862 163826 -1306
rect 164382 -1862 164414 -1306
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672618 167546 673174
rect 168102 672618 168134 673174
rect 167514 637174 168134 672618
rect 167514 636618 167546 637174
rect 168102 636618 168134 637174
rect 167514 601174 168134 636618
rect 167514 600618 167546 601174
rect 168102 600618 168134 601174
rect 167514 565174 168134 600618
rect 167514 564618 167546 565174
rect 168102 564618 168134 565174
rect 167514 529174 168134 564618
rect 167514 528618 167546 529174
rect 168102 528618 168134 529174
rect 167514 493174 168134 528618
rect 167514 492618 167546 493174
rect 168102 492618 168134 493174
rect 167514 457174 168134 492618
rect 167514 456618 167546 457174
rect 168102 456618 168134 457174
rect 167514 421174 168134 456618
rect 167514 420618 167546 421174
rect 168102 420618 168134 421174
rect 167514 385174 168134 420618
rect 167514 384618 167546 385174
rect 168102 384618 168134 385174
rect 167514 349174 168134 384618
rect 167514 348618 167546 349174
rect 168102 348618 168134 349174
rect 167514 313174 168134 348618
rect 167514 312618 167546 313174
rect 168102 312618 168134 313174
rect 167514 277174 168134 312618
rect 167514 276618 167546 277174
rect 168102 276618 168134 277174
rect 167514 241174 168134 276618
rect 167514 240618 167546 241174
rect 168102 240618 168134 241174
rect 167514 205174 168134 240618
rect 167514 204618 167546 205174
rect 168102 204618 168134 205174
rect 167514 169174 168134 204618
rect 167514 168618 167546 169174
rect 168102 168618 168134 169174
rect 167514 133174 168134 168618
rect 167514 132618 167546 133174
rect 168102 132618 168134 133174
rect 167514 97174 168134 132618
rect 167514 96618 167546 97174
rect 168102 96618 168134 97174
rect 167514 61174 168134 96618
rect 167514 60618 167546 61174
rect 168102 60618 168134 61174
rect 167514 25174 168134 60618
rect 167514 24618 167546 25174
rect 168102 24618 168134 25174
rect 167514 -3226 168134 24618
rect 167514 -3782 167546 -3226
rect 168102 -3782 168134 -3226
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676338 171266 676894
rect 171822 676338 171854 676894
rect 171234 640894 171854 676338
rect 171234 640338 171266 640894
rect 171822 640338 171854 640894
rect 171234 604894 171854 640338
rect 171234 604338 171266 604894
rect 171822 604338 171854 604894
rect 171234 568894 171854 604338
rect 171234 568338 171266 568894
rect 171822 568338 171854 568894
rect 171234 532894 171854 568338
rect 171234 532338 171266 532894
rect 171822 532338 171854 532894
rect 171234 496894 171854 532338
rect 171234 496338 171266 496894
rect 171822 496338 171854 496894
rect 171234 460894 171854 496338
rect 171234 460338 171266 460894
rect 171822 460338 171854 460894
rect 171234 424894 171854 460338
rect 171234 424338 171266 424894
rect 171822 424338 171854 424894
rect 171234 388894 171854 424338
rect 171234 388338 171266 388894
rect 171822 388338 171854 388894
rect 171234 352894 171854 388338
rect 171234 352338 171266 352894
rect 171822 352338 171854 352894
rect 171234 316894 171854 352338
rect 171234 316338 171266 316894
rect 171822 316338 171854 316894
rect 171234 280894 171854 316338
rect 171234 280338 171266 280894
rect 171822 280338 171854 280894
rect 171234 244894 171854 280338
rect 171234 244338 171266 244894
rect 171822 244338 171854 244894
rect 171234 208894 171854 244338
rect 171234 208338 171266 208894
rect 171822 208338 171854 208894
rect 171234 172894 171854 208338
rect 171234 172338 171266 172894
rect 171822 172338 171854 172894
rect 171234 136894 171854 172338
rect 171234 136338 171266 136894
rect 171822 136338 171854 136894
rect 171234 100894 171854 136338
rect 171234 100338 171266 100894
rect 171822 100338 171854 100894
rect 171234 64894 171854 100338
rect 171234 64338 171266 64894
rect 171822 64338 171854 64894
rect 171234 28894 171854 64338
rect 171234 28338 171266 28894
rect 171822 28338 171854 28894
rect 171234 -5146 171854 28338
rect 171234 -5702 171266 -5146
rect 171822 -5702 171854 -5146
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710042 192986 710598
rect 193542 710042 193574 710598
rect 189234 708678 189854 709670
rect 189234 708122 189266 708678
rect 189822 708122 189854 708678
rect 185514 706758 186134 707750
rect 185514 706202 185546 706758
rect 186102 706202 186134 706758
rect 174954 680058 174986 680614
rect 175542 680058 175574 680614
rect 174954 644614 175574 680058
rect 174954 644058 174986 644614
rect 175542 644058 175574 644614
rect 174954 608614 175574 644058
rect 174954 608058 174986 608614
rect 175542 608058 175574 608614
rect 174954 572614 175574 608058
rect 174954 572058 174986 572614
rect 175542 572058 175574 572614
rect 174954 536614 175574 572058
rect 174954 536058 174986 536614
rect 175542 536058 175574 536614
rect 174954 500614 175574 536058
rect 174954 500058 174986 500614
rect 175542 500058 175574 500614
rect 174954 464614 175574 500058
rect 174954 464058 174986 464614
rect 175542 464058 175574 464614
rect 174954 428614 175574 464058
rect 174954 428058 174986 428614
rect 175542 428058 175574 428614
rect 174954 392614 175574 428058
rect 174954 392058 174986 392614
rect 175542 392058 175574 392614
rect 174954 356614 175574 392058
rect 174954 356058 174986 356614
rect 175542 356058 175574 356614
rect 174954 320614 175574 356058
rect 174954 320058 174986 320614
rect 175542 320058 175574 320614
rect 174954 284614 175574 320058
rect 174954 284058 174986 284614
rect 175542 284058 175574 284614
rect 174954 248614 175574 284058
rect 174954 248058 174986 248614
rect 175542 248058 175574 248614
rect 174954 212614 175574 248058
rect 174954 212058 174986 212614
rect 175542 212058 175574 212614
rect 174954 176614 175574 212058
rect 174954 176058 174986 176614
rect 175542 176058 175574 176614
rect 174954 140614 175574 176058
rect 174954 140058 174986 140614
rect 175542 140058 175574 140614
rect 174954 104614 175574 140058
rect 174954 104058 174986 104614
rect 175542 104058 175574 104614
rect 174954 68614 175574 104058
rect 174954 68058 174986 68614
rect 175542 68058 175574 68614
rect 174954 32614 175574 68058
rect 174954 32058 174986 32614
rect 175542 32058 175574 32614
rect 156954 -6662 156986 -6106
rect 157542 -6662 157574 -6106
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704282 181826 704838
rect 182382 704282 182414 704838
rect 181794 687454 182414 704282
rect 181794 686898 181826 687454
rect 182382 686898 182414 687454
rect 181794 651454 182414 686898
rect 181794 650898 181826 651454
rect 182382 650898 182414 651454
rect 181794 615454 182414 650898
rect 181794 614898 181826 615454
rect 182382 614898 182414 615454
rect 181794 579454 182414 614898
rect 181794 578898 181826 579454
rect 182382 578898 182414 579454
rect 181794 543454 182414 578898
rect 181794 542898 181826 543454
rect 182382 542898 182414 543454
rect 181794 507454 182414 542898
rect 181794 506898 181826 507454
rect 182382 506898 182414 507454
rect 181794 471454 182414 506898
rect 181794 470898 181826 471454
rect 182382 470898 182414 471454
rect 181794 435454 182414 470898
rect 181794 434898 181826 435454
rect 182382 434898 182414 435454
rect 181794 399454 182414 434898
rect 181794 398898 181826 399454
rect 182382 398898 182414 399454
rect 181794 363454 182414 398898
rect 181794 362898 181826 363454
rect 182382 362898 182414 363454
rect 181794 327454 182414 362898
rect 181794 326898 181826 327454
rect 182382 326898 182414 327454
rect 181794 291454 182414 326898
rect 181794 290898 181826 291454
rect 182382 290898 182414 291454
rect 181794 255454 182414 290898
rect 181794 254898 181826 255454
rect 182382 254898 182414 255454
rect 181794 219454 182414 254898
rect 181794 218898 181826 219454
rect 182382 218898 182414 219454
rect 181794 183454 182414 218898
rect 181794 182898 181826 183454
rect 182382 182898 182414 183454
rect 181794 147454 182414 182898
rect 181794 146898 181826 147454
rect 182382 146898 182414 147454
rect 181794 111454 182414 146898
rect 181794 110898 181826 111454
rect 182382 110898 182414 111454
rect 181794 75454 182414 110898
rect 181794 74898 181826 75454
rect 182382 74898 182414 75454
rect 181794 39454 182414 74898
rect 181794 38898 181826 39454
rect 182382 38898 182414 39454
rect 181794 3454 182414 38898
rect 181794 2898 181826 3454
rect 182382 2898 182414 3454
rect 181794 -346 182414 2898
rect 181794 -902 181826 -346
rect 182382 -902 182414 -346
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690618 185546 691174
rect 186102 690618 186134 691174
rect 185514 655174 186134 690618
rect 185514 654618 185546 655174
rect 186102 654618 186134 655174
rect 185514 619174 186134 654618
rect 185514 618618 185546 619174
rect 186102 618618 186134 619174
rect 185514 583174 186134 618618
rect 185514 582618 185546 583174
rect 186102 582618 186134 583174
rect 185514 547174 186134 582618
rect 185514 546618 185546 547174
rect 186102 546618 186134 547174
rect 185514 511174 186134 546618
rect 185514 510618 185546 511174
rect 186102 510618 186134 511174
rect 185514 475174 186134 510618
rect 185514 474618 185546 475174
rect 186102 474618 186134 475174
rect 185514 439174 186134 474618
rect 185514 438618 185546 439174
rect 186102 438618 186134 439174
rect 185514 403174 186134 438618
rect 185514 402618 185546 403174
rect 186102 402618 186134 403174
rect 185514 367174 186134 402618
rect 185514 366618 185546 367174
rect 186102 366618 186134 367174
rect 185514 331174 186134 366618
rect 185514 330618 185546 331174
rect 186102 330618 186134 331174
rect 185514 295174 186134 330618
rect 185514 294618 185546 295174
rect 186102 294618 186134 295174
rect 185514 259174 186134 294618
rect 185514 258618 185546 259174
rect 186102 258618 186134 259174
rect 185514 223174 186134 258618
rect 185514 222618 185546 223174
rect 186102 222618 186134 223174
rect 185514 187174 186134 222618
rect 185514 186618 185546 187174
rect 186102 186618 186134 187174
rect 185514 151174 186134 186618
rect 185514 150618 185546 151174
rect 186102 150618 186134 151174
rect 185514 115174 186134 150618
rect 185514 114618 185546 115174
rect 186102 114618 186134 115174
rect 185514 79174 186134 114618
rect 185514 78618 185546 79174
rect 186102 78618 186134 79174
rect 185514 43174 186134 78618
rect 185514 42618 185546 43174
rect 186102 42618 186134 43174
rect 185514 7174 186134 42618
rect 185514 6618 185546 7174
rect 186102 6618 186134 7174
rect 185514 -2266 186134 6618
rect 185514 -2822 185546 -2266
rect 186102 -2822 186134 -2266
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694338 189266 694894
rect 189822 694338 189854 694894
rect 189234 658894 189854 694338
rect 189234 658338 189266 658894
rect 189822 658338 189854 658894
rect 189234 622894 189854 658338
rect 189234 622338 189266 622894
rect 189822 622338 189854 622894
rect 189234 586894 189854 622338
rect 189234 586338 189266 586894
rect 189822 586338 189854 586894
rect 189234 550894 189854 586338
rect 189234 550338 189266 550894
rect 189822 550338 189854 550894
rect 189234 514894 189854 550338
rect 189234 514338 189266 514894
rect 189822 514338 189854 514894
rect 189234 478894 189854 514338
rect 189234 478338 189266 478894
rect 189822 478338 189854 478894
rect 189234 442894 189854 478338
rect 189234 442338 189266 442894
rect 189822 442338 189854 442894
rect 189234 406894 189854 442338
rect 189234 406338 189266 406894
rect 189822 406338 189854 406894
rect 189234 370894 189854 406338
rect 189234 370338 189266 370894
rect 189822 370338 189854 370894
rect 189234 334894 189854 370338
rect 189234 334338 189266 334894
rect 189822 334338 189854 334894
rect 189234 298894 189854 334338
rect 189234 298338 189266 298894
rect 189822 298338 189854 298894
rect 189234 262894 189854 298338
rect 189234 262338 189266 262894
rect 189822 262338 189854 262894
rect 189234 226894 189854 262338
rect 189234 226338 189266 226894
rect 189822 226338 189854 226894
rect 189234 190894 189854 226338
rect 189234 190338 189266 190894
rect 189822 190338 189854 190894
rect 189234 154894 189854 190338
rect 189234 154338 189266 154894
rect 189822 154338 189854 154894
rect 189234 118894 189854 154338
rect 189234 118338 189266 118894
rect 189822 118338 189854 118894
rect 189234 82894 189854 118338
rect 189234 82338 189266 82894
rect 189822 82338 189854 82894
rect 189234 46894 189854 82338
rect 189234 46338 189266 46894
rect 189822 46338 189854 46894
rect 189234 10894 189854 46338
rect 189234 10338 189266 10894
rect 189822 10338 189854 10894
rect 189234 -4186 189854 10338
rect 189234 -4742 189266 -4186
rect 189822 -4742 189854 -4186
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711002 210986 711558
rect 211542 711002 211574 711558
rect 207234 709638 207854 709670
rect 207234 709082 207266 709638
rect 207822 709082 207854 709638
rect 203514 707718 204134 707750
rect 203514 707162 203546 707718
rect 204102 707162 204134 707718
rect 192954 698058 192986 698614
rect 193542 698058 193574 698614
rect 192954 662614 193574 698058
rect 192954 662058 192986 662614
rect 193542 662058 193574 662614
rect 192954 626614 193574 662058
rect 192954 626058 192986 626614
rect 193542 626058 193574 626614
rect 192954 590614 193574 626058
rect 192954 590058 192986 590614
rect 193542 590058 193574 590614
rect 192954 554614 193574 590058
rect 192954 554058 192986 554614
rect 193542 554058 193574 554614
rect 192954 518614 193574 554058
rect 192954 518058 192986 518614
rect 193542 518058 193574 518614
rect 192954 482614 193574 518058
rect 192954 482058 192986 482614
rect 193542 482058 193574 482614
rect 192954 446614 193574 482058
rect 192954 446058 192986 446614
rect 193542 446058 193574 446614
rect 192954 410614 193574 446058
rect 192954 410058 192986 410614
rect 193542 410058 193574 410614
rect 192954 374614 193574 410058
rect 192954 374058 192986 374614
rect 193542 374058 193574 374614
rect 192954 338614 193574 374058
rect 192954 338058 192986 338614
rect 193542 338058 193574 338614
rect 192954 302614 193574 338058
rect 192954 302058 192986 302614
rect 193542 302058 193574 302614
rect 192954 266614 193574 302058
rect 192954 266058 192986 266614
rect 193542 266058 193574 266614
rect 192954 230614 193574 266058
rect 192954 230058 192986 230614
rect 193542 230058 193574 230614
rect 192954 194614 193574 230058
rect 192954 194058 192986 194614
rect 193542 194058 193574 194614
rect 192954 158614 193574 194058
rect 192954 158058 192986 158614
rect 193542 158058 193574 158614
rect 192954 122614 193574 158058
rect 192954 122058 192986 122614
rect 193542 122058 193574 122614
rect 192954 86614 193574 122058
rect 192954 86058 192986 86614
rect 193542 86058 193574 86614
rect 192954 50614 193574 86058
rect 192954 50058 192986 50614
rect 193542 50058 193574 50614
rect 192954 14614 193574 50058
rect 192954 14058 192986 14614
rect 193542 14058 193574 14614
rect 174954 -7622 174986 -7066
rect 175542 -7622 175574 -7066
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705242 199826 705798
rect 200382 705242 200414 705798
rect 199794 669454 200414 705242
rect 199794 668898 199826 669454
rect 200382 668898 200414 669454
rect 199794 633454 200414 668898
rect 199794 632898 199826 633454
rect 200382 632898 200414 633454
rect 199794 597454 200414 632898
rect 199794 596898 199826 597454
rect 200382 596898 200414 597454
rect 199794 561454 200414 596898
rect 199794 560898 199826 561454
rect 200382 560898 200414 561454
rect 199794 525454 200414 560898
rect 199794 524898 199826 525454
rect 200382 524898 200414 525454
rect 199794 489454 200414 524898
rect 199794 488898 199826 489454
rect 200382 488898 200414 489454
rect 199794 453454 200414 488898
rect 199794 452898 199826 453454
rect 200382 452898 200414 453454
rect 199794 417454 200414 452898
rect 199794 416898 199826 417454
rect 200382 416898 200414 417454
rect 199794 381454 200414 416898
rect 199794 380898 199826 381454
rect 200382 380898 200414 381454
rect 199794 345454 200414 380898
rect 199794 344898 199826 345454
rect 200382 344898 200414 345454
rect 199794 309454 200414 344898
rect 199794 308898 199826 309454
rect 200382 308898 200414 309454
rect 199794 273454 200414 308898
rect 199794 272898 199826 273454
rect 200382 272898 200414 273454
rect 199794 237454 200414 272898
rect 199794 236898 199826 237454
rect 200382 236898 200414 237454
rect 199794 201454 200414 236898
rect 199794 200898 199826 201454
rect 200382 200898 200414 201454
rect 199794 165454 200414 200898
rect 199794 164898 199826 165454
rect 200382 164898 200414 165454
rect 199794 129454 200414 164898
rect 199794 128898 199826 129454
rect 200382 128898 200414 129454
rect 199794 93454 200414 128898
rect 199794 92898 199826 93454
rect 200382 92898 200414 93454
rect 199794 57454 200414 92898
rect 199794 56898 199826 57454
rect 200382 56898 200414 57454
rect 199794 21454 200414 56898
rect 199794 20898 199826 21454
rect 200382 20898 200414 21454
rect 199794 -1306 200414 20898
rect 199794 -1862 199826 -1306
rect 200382 -1862 200414 -1306
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672618 203546 673174
rect 204102 672618 204134 673174
rect 203514 637174 204134 672618
rect 203514 636618 203546 637174
rect 204102 636618 204134 637174
rect 203514 601174 204134 636618
rect 203514 600618 203546 601174
rect 204102 600618 204134 601174
rect 203514 565174 204134 600618
rect 203514 564618 203546 565174
rect 204102 564618 204134 565174
rect 203514 529174 204134 564618
rect 203514 528618 203546 529174
rect 204102 528618 204134 529174
rect 203514 493174 204134 528618
rect 203514 492618 203546 493174
rect 204102 492618 204134 493174
rect 203514 457174 204134 492618
rect 203514 456618 203546 457174
rect 204102 456618 204134 457174
rect 203514 421174 204134 456618
rect 203514 420618 203546 421174
rect 204102 420618 204134 421174
rect 203514 385174 204134 420618
rect 203514 384618 203546 385174
rect 204102 384618 204134 385174
rect 203514 349174 204134 384618
rect 203514 348618 203546 349174
rect 204102 348618 204134 349174
rect 203514 313174 204134 348618
rect 203514 312618 203546 313174
rect 204102 312618 204134 313174
rect 203514 277174 204134 312618
rect 203514 276618 203546 277174
rect 204102 276618 204134 277174
rect 203514 241174 204134 276618
rect 203514 240618 203546 241174
rect 204102 240618 204134 241174
rect 203514 205174 204134 240618
rect 203514 204618 203546 205174
rect 204102 204618 204134 205174
rect 203514 169174 204134 204618
rect 203514 168618 203546 169174
rect 204102 168618 204134 169174
rect 203514 133174 204134 168618
rect 203514 132618 203546 133174
rect 204102 132618 204134 133174
rect 203514 97174 204134 132618
rect 203514 96618 203546 97174
rect 204102 96618 204134 97174
rect 203514 61174 204134 96618
rect 203514 60618 203546 61174
rect 204102 60618 204134 61174
rect 203514 25174 204134 60618
rect 203514 24618 203546 25174
rect 204102 24618 204134 25174
rect 203514 -3226 204134 24618
rect 203514 -3782 203546 -3226
rect 204102 -3782 204134 -3226
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676338 207266 676894
rect 207822 676338 207854 676894
rect 207234 640894 207854 676338
rect 207234 640338 207266 640894
rect 207822 640338 207854 640894
rect 207234 604894 207854 640338
rect 207234 604338 207266 604894
rect 207822 604338 207854 604894
rect 207234 568894 207854 604338
rect 207234 568338 207266 568894
rect 207822 568338 207854 568894
rect 207234 532894 207854 568338
rect 207234 532338 207266 532894
rect 207822 532338 207854 532894
rect 207234 496894 207854 532338
rect 207234 496338 207266 496894
rect 207822 496338 207854 496894
rect 207234 460894 207854 496338
rect 207234 460338 207266 460894
rect 207822 460338 207854 460894
rect 207234 424894 207854 460338
rect 207234 424338 207266 424894
rect 207822 424338 207854 424894
rect 207234 388894 207854 424338
rect 207234 388338 207266 388894
rect 207822 388338 207854 388894
rect 207234 352894 207854 388338
rect 207234 352338 207266 352894
rect 207822 352338 207854 352894
rect 207234 316894 207854 352338
rect 207234 316338 207266 316894
rect 207822 316338 207854 316894
rect 207234 280894 207854 316338
rect 207234 280338 207266 280894
rect 207822 280338 207854 280894
rect 207234 244894 207854 280338
rect 207234 244338 207266 244894
rect 207822 244338 207854 244894
rect 207234 208894 207854 244338
rect 207234 208338 207266 208894
rect 207822 208338 207854 208894
rect 207234 172894 207854 208338
rect 207234 172338 207266 172894
rect 207822 172338 207854 172894
rect 207234 136894 207854 172338
rect 207234 136338 207266 136894
rect 207822 136338 207854 136894
rect 207234 100894 207854 136338
rect 207234 100338 207266 100894
rect 207822 100338 207854 100894
rect 207234 64894 207854 100338
rect 207234 64338 207266 64894
rect 207822 64338 207854 64894
rect 207234 28894 207854 64338
rect 207234 28338 207266 28894
rect 207822 28338 207854 28894
rect 207234 -5146 207854 28338
rect 207234 -5702 207266 -5146
rect 207822 -5702 207854 -5146
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710042 228986 710598
rect 229542 710042 229574 710598
rect 225234 708678 225854 709670
rect 225234 708122 225266 708678
rect 225822 708122 225854 708678
rect 221514 706758 222134 707750
rect 221514 706202 221546 706758
rect 222102 706202 222134 706758
rect 210954 680058 210986 680614
rect 211542 680058 211574 680614
rect 210954 644614 211574 680058
rect 210954 644058 210986 644614
rect 211542 644058 211574 644614
rect 210954 608614 211574 644058
rect 210954 608058 210986 608614
rect 211542 608058 211574 608614
rect 210954 572614 211574 608058
rect 210954 572058 210986 572614
rect 211542 572058 211574 572614
rect 210954 536614 211574 572058
rect 210954 536058 210986 536614
rect 211542 536058 211574 536614
rect 210954 500614 211574 536058
rect 210954 500058 210986 500614
rect 211542 500058 211574 500614
rect 210954 464614 211574 500058
rect 210954 464058 210986 464614
rect 211542 464058 211574 464614
rect 210954 428614 211574 464058
rect 210954 428058 210986 428614
rect 211542 428058 211574 428614
rect 210954 392614 211574 428058
rect 210954 392058 210986 392614
rect 211542 392058 211574 392614
rect 210954 356614 211574 392058
rect 210954 356058 210986 356614
rect 211542 356058 211574 356614
rect 210954 320614 211574 356058
rect 210954 320058 210986 320614
rect 211542 320058 211574 320614
rect 210954 284614 211574 320058
rect 210954 284058 210986 284614
rect 211542 284058 211574 284614
rect 210954 248614 211574 284058
rect 210954 248058 210986 248614
rect 211542 248058 211574 248614
rect 210954 212614 211574 248058
rect 210954 212058 210986 212614
rect 211542 212058 211574 212614
rect 210954 176614 211574 212058
rect 210954 176058 210986 176614
rect 211542 176058 211574 176614
rect 210954 140614 211574 176058
rect 210954 140058 210986 140614
rect 211542 140058 211574 140614
rect 210954 104614 211574 140058
rect 210954 104058 210986 104614
rect 211542 104058 211574 104614
rect 210954 68614 211574 104058
rect 210954 68058 210986 68614
rect 211542 68058 211574 68614
rect 210954 32614 211574 68058
rect 210954 32058 210986 32614
rect 211542 32058 211574 32614
rect 192954 -6662 192986 -6106
rect 193542 -6662 193574 -6106
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704282 217826 704838
rect 218382 704282 218414 704838
rect 217794 687454 218414 704282
rect 217794 686898 217826 687454
rect 218382 686898 218414 687454
rect 217794 651454 218414 686898
rect 217794 650898 217826 651454
rect 218382 650898 218414 651454
rect 217794 615454 218414 650898
rect 217794 614898 217826 615454
rect 218382 614898 218414 615454
rect 217794 579454 218414 614898
rect 217794 578898 217826 579454
rect 218382 578898 218414 579454
rect 217794 543454 218414 578898
rect 217794 542898 217826 543454
rect 218382 542898 218414 543454
rect 217794 507454 218414 542898
rect 217794 506898 217826 507454
rect 218382 506898 218414 507454
rect 217794 471454 218414 506898
rect 217794 470898 217826 471454
rect 218382 470898 218414 471454
rect 217794 435454 218414 470898
rect 217794 434898 217826 435454
rect 218382 434898 218414 435454
rect 217794 399454 218414 434898
rect 217794 398898 217826 399454
rect 218382 398898 218414 399454
rect 217794 363454 218414 398898
rect 217794 362898 217826 363454
rect 218382 362898 218414 363454
rect 217794 327454 218414 362898
rect 217794 326898 217826 327454
rect 218382 326898 218414 327454
rect 217794 291454 218414 326898
rect 217794 290898 217826 291454
rect 218382 290898 218414 291454
rect 217794 255454 218414 290898
rect 217794 254898 217826 255454
rect 218382 254898 218414 255454
rect 217794 219454 218414 254898
rect 217794 218898 217826 219454
rect 218382 218898 218414 219454
rect 217794 183454 218414 218898
rect 217794 182898 217826 183454
rect 218382 182898 218414 183454
rect 217794 147454 218414 182898
rect 217794 146898 217826 147454
rect 218382 146898 218414 147454
rect 217794 111454 218414 146898
rect 217794 110898 217826 111454
rect 218382 110898 218414 111454
rect 217794 75454 218414 110898
rect 217794 74898 217826 75454
rect 218382 74898 218414 75454
rect 217794 39454 218414 74898
rect 217794 38898 217826 39454
rect 218382 38898 218414 39454
rect 217794 3454 218414 38898
rect 217794 2898 217826 3454
rect 218382 2898 218414 3454
rect 217794 -346 218414 2898
rect 217794 -902 217826 -346
rect 218382 -902 218414 -346
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690618 221546 691174
rect 222102 690618 222134 691174
rect 221514 655174 222134 690618
rect 221514 654618 221546 655174
rect 222102 654618 222134 655174
rect 221514 619174 222134 654618
rect 221514 618618 221546 619174
rect 222102 618618 222134 619174
rect 221514 583174 222134 618618
rect 221514 582618 221546 583174
rect 222102 582618 222134 583174
rect 221514 547174 222134 582618
rect 221514 546618 221546 547174
rect 222102 546618 222134 547174
rect 221514 511174 222134 546618
rect 221514 510618 221546 511174
rect 222102 510618 222134 511174
rect 221514 475174 222134 510618
rect 221514 474618 221546 475174
rect 222102 474618 222134 475174
rect 221514 439174 222134 474618
rect 221514 438618 221546 439174
rect 222102 438618 222134 439174
rect 221514 403174 222134 438618
rect 221514 402618 221546 403174
rect 222102 402618 222134 403174
rect 221514 367174 222134 402618
rect 221514 366618 221546 367174
rect 222102 366618 222134 367174
rect 221514 331174 222134 366618
rect 221514 330618 221546 331174
rect 222102 330618 222134 331174
rect 221514 295174 222134 330618
rect 221514 294618 221546 295174
rect 222102 294618 222134 295174
rect 221514 259174 222134 294618
rect 221514 258618 221546 259174
rect 222102 258618 222134 259174
rect 221514 223174 222134 258618
rect 221514 222618 221546 223174
rect 222102 222618 222134 223174
rect 221514 187174 222134 222618
rect 221514 186618 221546 187174
rect 222102 186618 222134 187174
rect 221514 151174 222134 186618
rect 221514 150618 221546 151174
rect 222102 150618 222134 151174
rect 221514 115174 222134 150618
rect 221514 114618 221546 115174
rect 222102 114618 222134 115174
rect 221514 79174 222134 114618
rect 221514 78618 221546 79174
rect 222102 78618 222134 79174
rect 221514 43174 222134 78618
rect 221514 42618 221546 43174
rect 222102 42618 222134 43174
rect 221514 7174 222134 42618
rect 221514 6618 221546 7174
rect 222102 6618 222134 7174
rect 221514 -2266 222134 6618
rect 221514 -2822 221546 -2266
rect 222102 -2822 222134 -2266
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694338 225266 694894
rect 225822 694338 225854 694894
rect 225234 658894 225854 694338
rect 225234 658338 225266 658894
rect 225822 658338 225854 658894
rect 225234 622894 225854 658338
rect 225234 622338 225266 622894
rect 225822 622338 225854 622894
rect 225234 586894 225854 622338
rect 225234 586338 225266 586894
rect 225822 586338 225854 586894
rect 225234 550894 225854 586338
rect 225234 550338 225266 550894
rect 225822 550338 225854 550894
rect 225234 514894 225854 550338
rect 225234 514338 225266 514894
rect 225822 514338 225854 514894
rect 225234 478894 225854 514338
rect 225234 478338 225266 478894
rect 225822 478338 225854 478894
rect 225234 442894 225854 478338
rect 225234 442338 225266 442894
rect 225822 442338 225854 442894
rect 225234 406894 225854 442338
rect 225234 406338 225266 406894
rect 225822 406338 225854 406894
rect 225234 370894 225854 406338
rect 225234 370338 225266 370894
rect 225822 370338 225854 370894
rect 225234 334894 225854 370338
rect 225234 334338 225266 334894
rect 225822 334338 225854 334894
rect 225234 298894 225854 334338
rect 225234 298338 225266 298894
rect 225822 298338 225854 298894
rect 225234 262894 225854 298338
rect 225234 262338 225266 262894
rect 225822 262338 225854 262894
rect 225234 226894 225854 262338
rect 225234 226338 225266 226894
rect 225822 226338 225854 226894
rect 225234 190894 225854 226338
rect 225234 190338 225266 190894
rect 225822 190338 225854 190894
rect 225234 154894 225854 190338
rect 225234 154338 225266 154894
rect 225822 154338 225854 154894
rect 225234 118894 225854 154338
rect 225234 118338 225266 118894
rect 225822 118338 225854 118894
rect 225234 82894 225854 118338
rect 225234 82338 225266 82894
rect 225822 82338 225854 82894
rect 225234 46894 225854 82338
rect 225234 46338 225266 46894
rect 225822 46338 225854 46894
rect 225234 10894 225854 46338
rect 225234 10338 225266 10894
rect 225822 10338 225854 10894
rect 225234 -4186 225854 10338
rect 225234 -4742 225266 -4186
rect 225822 -4742 225854 -4186
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711002 246986 711558
rect 247542 711002 247574 711558
rect 243234 709638 243854 709670
rect 243234 709082 243266 709638
rect 243822 709082 243854 709638
rect 239514 707718 240134 707750
rect 239514 707162 239546 707718
rect 240102 707162 240134 707718
rect 228954 698058 228986 698614
rect 229542 698058 229574 698614
rect 228954 662614 229574 698058
rect 228954 662058 228986 662614
rect 229542 662058 229574 662614
rect 228954 626614 229574 662058
rect 228954 626058 228986 626614
rect 229542 626058 229574 626614
rect 228954 590614 229574 626058
rect 228954 590058 228986 590614
rect 229542 590058 229574 590614
rect 228954 554614 229574 590058
rect 228954 554058 228986 554614
rect 229542 554058 229574 554614
rect 228954 518614 229574 554058
rect 228954 518058 228986 518614
rect 229542 518058 229574 518614
rect 228954 482614 229574 518058
rect 235794 705798 236414 705830
rect 235794 705242 235826 705798
rect 236382 705242 236414 705798
rect 235794 669454 236414 705242
rect 235794 668898 235826 669454
rect 236382 668898 236414 669454
rect 235794 633454 236414 668898
rect 235794 632898 235826 633454
rect 236382 632898 236414 633454
rect 235794 597454 236414 632898
rect 235794 596898 235826 597454
rect 236382 596898 236414 597454
rect 235794 561454 236414 596898
rect 235794 560898 235826 561454
rect 236382 560898 236414 561454
rect 235794 525454 236414 560898
rect 235794 524898 235826 525454
rect 236382 524898 236414 525454
rect 235794 500000 236414 524898
rect 239514 673174 240134 707162
rect 239514 672618 239546 673174
rect 240102 672618 240134 673174
rect 239514 637174 240134 672618
rect 239514 636618 239546 637174
rect 240102 636618 240134 637174
rect 239514 601174 240134 636618
rect 239514 600618 239546 601174
rect 240102 600618 240134 601174
rect 239514 565174 240134 600618
rect 239514 564618 239546 565174
rect 240102 564618 240134 565174
rect 239514 529174 240134 564618
rect 239514 528618 239546 529174
rect 240102 528618 240134 529174
rect 236683 500308 236749 500309
rect 236683 500244 236684 500308
rect 236748 500244 236749 500308
rect 236683 500243 236749 500244
rect 236499 500172 236565 500173
rect 236499 500108 236500 500172
rect 236564 500108 236565 500172
rect 236499 500107 236565 500108
rect 233739 498676 233805 498677
rect 233739 498612 233740 498676
rect 233804 498612 233805 498676
rect 233739 498611 233805 498612
rect 228954 482058 228986 482614
rect 229542 482058 229574 482614
rect 228954 446614 229574 482058
rect 228954 446058 228986 446614
rect 229542 446058 229574 446614
rect 228954 410614 229574 446058
rect 228954 410058 228986 410614
rect 229542 410058 229574 410614
rect 228954 374614 229574 410058
rect 228954 374058 228986 374614
rect 229542 374058 229574 374614
rect 228954 338614 229574 374058
rect 228954 338058 228986 338614
rect 229542 338058 229574 338614
rect 228954 302614 229574 338058
rect 228954 302058 228986 302614
rect 229542 302058 229574 302614
rect 228954 266614 229574 302058
rect 228954 266058 228986 266614
rect 229542 266058 229574 266614
rect 228954 230614 229574 266058
rect 228954 230058 228986 230614
rect 229542 230058 229574 230614
rect 228954 194614 229574 230058
rect 228954 194058 228986 194614
rect 229542 194058 229574 194614
rect 228954 158614 229574 194058
rect 228954 158058 228986 158614
rect 229542 158058 229574 158614
rect 228954 122614 229574 158058
rect 228954 122058 228986 122614
rect 229542 122058 229574 122614
rect 228954 86614 229574 122058
rect 228954 86058 228986 86614
rect 229542 86058 229574 86614
rect 228954 50614 229574 86058
rect 233742 84285 233802 498611
rect 235794 309454 236414 336000
rect 235794 308898 235826 309454
rect 236382 308898 236414 309454
rect 235794 273454 236414 308898
rect 235794 272898 235826 273454
rect 236382 272898 236414 273454
rect 235794 237454 236414 272898
rect 236502 266389 236562 500107
rect 236686 318885 236746 500243
rect 239514 500000 240134 528618
rect 243234 676894 243854 709082
rect 243234 676338 243266 676894
rect 243822 676338 243854 676894
rect 243234 640894 243854 676338
rect 243234 640338 243266 640894
rect 243822 640338 243854 640894
rect 243234 604894 243854 640338
rect 243234 604338 243266 604894
rect 243822 604338 243854 604894
rect 243234 568894 243854 604338
rect 243234 568338 243266 568894
rect 243822 568338 243854 568894
rect 243234 532894 243854 568338
rect 243234 532338 243266 532894
rect 243822 532338 243854 532894
rect 243234 500000 243854 532338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710042 264986 710598
rect 265542 710042 265574 710598
rect 261234 708678 261854 709670
rect 261234 708122 261266 708678
rect 261822 708122 261854 708678
rect 257514 706758 258134 707750
rect 257514 706202 257546 706758
rect 258102 706202 258134 706758
rect 246954 680058 246986 680614
rect 247542 680058 247574 680614
rect 246954 644614 247574 680058
rect 246954 644058 246986 644614
rect 247542 644058 247574 644614
rect 246954 608614 247574 644058
rect 246954 608058 246986 608614
rect 247542 608058 247574 608614
rect 246954 572614 247574 608058
rect 246954 572058 246986 572614
rect 247542 572058 247574 572614
rect 246954 536614 247574 572058
rect 246954 536058 246986 536614
rect 247542 536058 247574 536614
rect 246954 500614 247574 536058
rect 246954 500058 246986 500614
rect 247542 500058 247574 500614
rect 246954 500000 247574 500058
rect 253794 704838 254414 705830
rect 253794 704282 253826 704838
rect 254382 704282 254414 704838
rect 253794 687454 254414 704282
rect 253794 686898 253826 687454
rect 254382 686898 254414 687454
rect 253794 651454 254414 686898
rect 253794 650898 253826 651454
rect 254382 650898 254414 651454
rect 253794 615454 254414 650898
rect 253794 614898 253826 615454
rect 254382 614898 254414 615454
rect 253794 579454 254414 614898
rect 253794 578898 253826 579454
rect 254382 578898 254414 579454
rect 253794 543454 254414 578898
rect 253794 542898 253826 543454
rect 254382 542898 254414 543454
rect 253794 507454 254414 542898
rect 253794 506898 253826 507454
rect 254382 506898 254414 507454
rect 253794 500000 254414 506898
rect 257514 691174 258134 706202
rect 257514 690618 257546 691174
rect 258102 690618 258134 691174
rect 257514 655174 258134 690618
rect 257514 654618 257546 655174
rect 258102 654618 258134 655174
rect 257514 619174 258134 654618
rect 257514 618618 257546 619174
rect 258102 618618 258134 619174
rect 257514 583174 258134 618618
rect 257514 582618 257546 583174
rect 258102 582618 258134 583174
rect 257514 547174 258134 582618
rect 257514 546618 257546 547174
rect 258102 546618 258134 547174
rect 257514 511174 258134 546618
rect 257514 510618 257546 511174
rect 258102 510618 258134 511174
rect 257514 500000 258134 510618
rect 261234 694894 261854 708122
rect 261234 694338 261266 694894
rect 261822 694338 261854 694894
rect 261234 658894 261854 694338
rect 261234 658338 261266 658894
rect 261822 658338 261854 658894
rect 261234 622894 261854 658338
rect 261234 622338 261266 622894
rect 261822 622338 261854 622894
rect 261234 586894 261854 622338
rect 261234 586338 261266 586894
rect 261822 586338 261854 586894
rect 261234 550894 261854 586338
rect 261234 550338 261266 550894
rect 261822 550338 261854 550894
rect 261234 514894 261854 550338
rect 261234 514338 261266 514894
rect 261822 514338 261854 514894
rect 261234 500000 261854 514338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711002 282986 711558
rect 283542 711002 283574 711558
rect 279234 709638 279854 709670
rect 279234 709082 279266 709638
rect 279822 709082 279854 709638
rect 275514 707718 276134 707750
rect 275514 707162 275546 707718
rect 276102 707162 276134 707718
rect 264954 698058 264986 698614
rect 265542 698058 265574 698614
rect 264954 662614 265574 698058
rect 264954 662058 264986 662614
rect 265542 662058 265574 662614
rect 264954 626614 265574 662058
rect 264954 626058 264986 626614
rect 265542 626058 265574 626614
rect 264954 590614 265574 626058
rect 264954 590058 264986 590614
rect 265542 590058 265574 590614
rect 264954 554614 265574 590058
rect 264954 554058 264986 554614
rect 265542 554058 265574 554614
rect 264954 518614 265574 554058
rect 264954 518058 264986 518614
rect 265542 518058 265574 518614
rect 264954 500000 265574 518058
rect 271794 705798 272414 705830
rect 271794 705242 271826 705798
rect 272382 705242 272414 705798
rect 271794 669454 272414 705242
rect 271794 668898 271826 669454
rect 272382 668898 272414 669454
rect 271794 633454 272414 668898
rect 271794 632898 271826 633454
rect 272382 632898 272414 633454
rect 271794 597454 272414 632898
rect 271794 596898 271826 597454
rect 272382 596898 272414 597454
rect 271794 561454 272414 596898
rect 271794 560898 271826 561454
rect 272382 560898 272414 561454
rect 271794 525454 272414 560898
rect 271794 524898 271826 525454
rect 272382 524898 272414 525454
rect 271794 500000 272414 524898
rect 275514 673174 276134 707162
rect 275514 672618 275546 673174
rect 276102 672618 276134 673174
rect 275514 637174 276134 672618
rect 275514 636618 275546 637174
rect 276102 636618 276134 637174
rect 275514 601174 276134 636618
rect 275514 600618 275546 601174
rect 276102 600618 276134 601174
rect 275514 565174 276134 600618
rect 275514 564618 275546 565174
rect 276102 564618 276134 565174
rect 275514 529174 276134 564618
rect 275514 528618 275546 529174
rect 276102 528618 276134 529174
rect 275514 500000 276134 528618
rect 279234 676894 279854 709082
rect 279234 676338 279266 676894
rect 279822 676338 279854 676894
rect 279234 640894 279854 676338
rect 279234 640338 279266 640894
rect 279822 640338 279854 640894
rect 279234 604894 279854 640338
rect 279234 604338 279266 604894
rect 279822 604338 279854 604894
rect 279234 568894 279854 604338
rect 279234 568338 279266 568894
rect 279822 568338 279854 568894
rect 279234 532894 279854 568338
rect 279234 532338 279266 532894
rect 279822 532338 279854 532894
rect 279234 500000 279854 532338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710042 300986 710598
rect 301542 710042 301574 710598
rect 297234 708678 297854 709670
rect 297234 708122 297266 708678
rect 297822 708122 297854 708678
rect 293514 706758 294134 707750
rect 293514 706202 293546 706758
rect 294102 706202 294134 706758
rect 282954 680058 282986 680614
rect 283542 680058 283574 680614
rect 282954 644614 283574 680058
rect 282954 644058 282986 644614
rect 283542 644058 283574 644614
rect 282954 608614 283574 644058
rect 282954 608058 282986 608614
rect 283542 608058 283574 608614
rect 282954 572614 283574 608058
rect 282954 572058 282986 572614
rect 283542 572058 283574 572614
rect 282954 536614 283574 572058
rect 282954 536058 282986 536614
rect 283542 536058 283574 536614
rect 282954 500614 283574 536058
rect 282954 500058 282986 500614
rect 283542 500058 283574 500614
rect 282954 500000 283574 500058
rect 289794 704838 290414 705830
rect 289794 704282 289826 704838
rect 290382 704282 290414 704838
rect 289794 687454 290414 704282
rect 289794 686898 289826 687454
rect 290382 686898 290414 687454
rect 289794 651454 290414 686898
rect 289794 650898 289826 651454
rect 290382 650898 290414 651454
rect 289794 615454 290414 650898
rect 289794 614898 289826 615454
rect 290382 614898 290414 615454
rect 289794 579454 290414 614898
rect 289794 578898 289826 579454
rect 290382 578898 290414 579454
rect 289794 543454 290414 578898
rect 289794 542898 289826 543454
rect 290382 542898 290414 543454
rect 289794 507454 290414 542898
rect 289794 506898 289826 507454
rect 290382 506898 290414 507454
rect 289794 500000 290414 506898
rect 293514 691174 294134 706202
rect 293514 690618 293546 691174
rect 294102 690618 294134 691174
rect 293514 655174 294134 690618
rect 293514 654618 293546 655174
rect 294102 654618 294134 655174
rect 293514 619174 294134 654618
rect 293514 618618 293546 619174
rect 294102 618618 294134 619174
rect 293514 583174 294134 618618
rect 293514 582618 293546 583174
rect 294102 582618 294134 583174
rect 293514 547174 294134 582618
rect 293514 546618 293546 547174
rect 294102 546618 294134 547174
rect 293514 511174 294134 546618
rect 293514 510618 293546 511174
rect 294102 510618 294134 511174
rect 293514 500000 294134 510618
rect 297234 694894 297854 708122
rect 297234 694338 297266 694894
rect 297822 694338 297854 694894
rect 297234 658894 297854 694338
rect 297234 658338 297266 658894
rect 297822 658338 297854 658894
rect 297234 622894 297854 658338
rect 297234 622338 297266 622894
rect 297822 622338 297854 622894
rect 297234 586894 297854 622338
rect 297234 586338 297266 586894
rect 297822 586338 297854 586894
rect 297234 550894 297854 586338
rect 297234 550338 297266 550894
rect 297822 550338 297854 550894
rect 297234 514894 297854 550338
rect 297234 514338 297266 514894
rect 297822 514338 297854 514894
rect 297234 500000 297854 514338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711002 318986 711558
rect 319542 711002 319574 711558
rect 315234 709638 315854 709670
rect 315234 709082 315266 709638
rect 315822 709082 315854 709638
rect 311514 707718 312134 707750
rect 311514 707162 311546 707718
rect 312102 707162 312134 707718
rect 300954 698058 300986 698614
rect 301542 698058 301574 698614
rect 300954 662614 301574 698058
rect 300954 662058 300986 662614
rect 301542 662058 301574 662614
rect 300954 626614 301574 662058
rect 300954 626058 300986 626614
rect 301542 626058 301574 626614
rect 300954 590614 301574 626058
rect 300954 590058 300986 590614
rect 301542 590058 301574 590614
rect 300954 554614 301574 590058
rect 300954 554058 300986 554614
rect 301542 554058 301574 554614
rect 300954 518614 301574 554058
rect 300954 518058 300986 518614
rect 301542 518058 301574 518614
rect 300954 500000 301574 518058
rect 307794 705798 308414 705830
rect 307794 705242 307826 705798
rect 308382 705242 308414 705798
rect 307794 669454 308414 705242
rect 307794 668898 307826 669454
rect 308382 668898 308414 669454
rect 307794 633454 308414 668898
rect 307794 632898 307826 633454
rect 308382 632898 308414 633454
rect 307794 597454 308414 632898
rect 307794 596898 307826 597454
rect 308382 596898 308414 597454
rect 307794 561454 308414 596898
rect 307794 560898 307826 561454
rect 308382 560898 308414 561454
rect 307794 525454 308414 560898
rect 307794 524898 307826 525454
rect 308382 524898 308414 525454
rect 307794 500000 308414 524898
rect 311514 673174 312134 707162
rect 311514 672618 311546 673174
rect 312102 672618 312134 673174
rect 311514 637174 312134 672618
rect 311514 636618 311546 637174
rect 312102 636618 312134 637174
rect 311514 601174 312134 636618
rect 311514 600618 311546 601174
rect 312102 600618 312134 601174
rect 311514 565174 312134 600618
rect 311514 564618 311546 565174
rect 312102 564618 312134 565174
rect 311514 529174 312134 564618
rect 311514 528618 311546 529174
rect 312102 528618 312134 529174
rect 311514 500000 312134 528618
rect 315234 676894 315854 709082
rect 315234 676338 315266 676894
rect 315822 676338 315854 676894
rect 315234 640894 315854 676338
rect 315234 640338 315266 640894
rect 315822 640338 315854 640894
rect 315234 604894 315854 640338
rect 315234 604338 315266 604894
rect 315822 604338 315854 604894
rect 315234 568894 315854 604338
rect 315234 568338 315266 568894
rect 315822 568338 315854 568894
rect 315234 532894 315854 568338
rect 315234 532338 315266 532894
rect 315822 532338 315854 532894
rect 315234 500000 315854 532338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710042 336986 710598
rect 337542 710042 337574 710598
rect 333234 708678 333854 709670
rect 333234 708122 333266 708678
rect 333822 708122 333854 708678
rect 329514 706758 330134 707750
rect 329514 706202 329546 706758
rect 330102 706202 330134 706758
rect 318954 680058 318986 680614
rect 319542 680058 319574 680614
rect 318954 644614 319574 680058
rect 318954 644058 318986 644614
rect 319542 644058 319574 644614
rect 318954 608614 319574 644058
rect 318954 608058 318986 608614
rect 319542 608058 319574 608614
rect 318954 572614 319574 608058
rect 318954 572058 318986 572614
rect 319542 572058 319574 572614
rect 318954 536614 319574 572058
rect 318954 536058 318986 536614
rect 319542 536058 319574 536614
rect 318954 500614 319574 536058
rect 318954 500058 318986 500614
rect 319542 500058 319574 500614
rect 318954 500000 319574 500058
rect 325794 704838 326414 705830
rect 325794 704282 325826 704838
rect 326382 704282 326414 704838
rect 325794 687454 326414 704282
rect 325794 686898 325826 687454
rect 326382 686898 326414 687454
rect 325794 651454 326414 686898
rect 325794 650898 325826 651454
rect 326382 650898 326414 651454
rect 325794 615454 326414 650898
rect 325794 614898 325826 615454
rect 326382 614898 326414 615454
rect 325794 579454 326414 614898
rect 325794 578898 325826 579454
rect 326382 578898 326414 579454
rect 325794 543454 326414 578898
rect 325794 542898 325826 543454
rect 326382 542898 326414 543454
rect 325794 507454 326414 542898
rect 325794 506898 325826 507454
rect 326382 506898 326414 507454
rect 325794 500000 326414 506898
rect 329514 691174 330134 706202
rect 329514 690618 329546 691174
rect 330102 690618 330134 691174
rect 329514 655174 330134 690618
rect 329514 654618 329546 655174
rect 330102 654618 330134 655174
rect 329514 619174 330134 654618
rect 329514 618618 329546 619174
rect 330102 618618 330134 619174
rect 329514 583174 330134 618618
rect 329514 582618 329546 583174
rect 330102 582618 330134 583174
rect 329514 547174 330134 582618
rect 329514 546618 329546 547174
rect 330102 546618 330134 547174
rect 329514 511174 330134 546618
rect 329514 510618 329546 511174
rect 330102 510618 330134 511174
rect 329514 500000 330134 510618
rect 333234 694894 333854 708122
rect 333234 694338 333266 694894
rect 333822 694338 333854 694894
rect 333234 658894 333854 694338
rect 333234 658338 333266 658894
rect 333822 658338 333854 658894
rect 333234 622894 333854 658338
rect 333234 622338 333266 622894
rect 333822 622338 333854 622894
rect 333234 586894 333854 622338
rect 333234 586338 333266 586894
rect 333822 586338 333854 586894
rect 333234 550894 333854 586338
rect 333234 550338 333266 550894
rect 333822 550338 333854 550894
rect 333234 514894 333854 550338
rect 333234 514338 333266 514894
rect 333822 514338 333854 514894
rect 333234 500000 333854 514338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711002 354986 711558
rect 355542 711002 355574 711558
rect 351234 709638 351854 709670
rect 351234 709082 351266 709638
rect 351822 709082 351854 709638
rect 347514 707718 348134 707750
rect 347514 707162 347546 707718
rect 348102 707162 348134 707718
rect 336954 698058 336986 698614
rect 337542 698058 337574 698614
rect 336954 662614 337574 698058
rect 336954 662058 336986 662614
rect 337542 662058 337574 662614
rect 336954 626614 337574 662058
rect 336954 626058 336986 626614
rect 337542 626058 337574 626614
rect 336954 590614 337574 626058
rect 336954 590058 336986 590614
rect 337542 590058 337574 590614
rect 336954 554614 337574 590058
rect 336954 554058 336986 554614
rect 337542 554058 337574 554614
rect 336954 518614 337574 554058
rect 336954 518058 336986 518614
rect 337542 518058 337574 518614
rect 336954 500000 337574 518058
rect 343794 705798 344414 705830
rect 343794 705242 343826 705798
rect 344382 705242 344414 705798
rect 343794 669454 344414 705242
rect 343794 668898 343826 669454
rect 344382 668898 344414 669454
rect 343794 633454 344414 668898
rect 343794 632898 343826 633454
rect 344382 632898 344414 633454
rect 343794 597454 344414 632898
rect 343794 596898 343826 597454
rect 344382 596898 344414 597454
rect 343794 561454 344414 596898
rect 343794 560898 343826 561454
rect 344382 560898 344414 561454
rect 343794 525454 344414 560898
rect 343794 524898 343826 525454
rect 344382 524898 344414 525454
rect 343794 500000 344414 524898
rect 347514 673174 348134 707162
rect 347514 672618 347546 673174
rect 348102 672618 348134 673174
rect 347514 637174 348134 672618
rect 347514 636618 347546 637174
rect 348102 636618 348134 637174
rect 347514 601174 348134 636618
rect 347514 600618 347546 601174
rect 348102 600618 348134 601174
rect 347514 565174 348134 600618
rect 347514 564618 347546 565174
rect 348102 564618 348134 565174
rect 347514 529174 348134 564618
rect 347514 528618 347546 529174
rect 348102 528618 348134 529174
rect 347514 500000 348134 528618
rect 351234 676894 351854 709082
rect 351234 676338 351266 676894
rect 351822 676338 351854 676894
rect 351234 640894 351854 676338
rect 351234 640338 351266 640894
rect 351822 640338 351854 640894
rect 351234 604894 351854 640338
rect 351234 604338 351266 604894
rect 351822 604338 351854 604894
rect 351234 568894 351854 604338
rect 351234 568338 351266 568894
rect 351822 568338 351854 568894
rect 351234 532894 351854 568338
rect 351234 532338 351266 532894
rect 351822 532338 351854 532894
rect 351234 500000 351854 532338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710042 372986 710598
rect 373542 710042 373574 710598
rect 369234 708678 369854 709670
rect 369234 708122 369266 708678
rect 369822 708122 369854 708678
rect 365514 706758 366134 707750
rect 365514 706202 365546 706758
rect 366102 706202 366134 706758
rect 354954 680058 354986 680614
rect 355542 680058 355574 680614
rect 354954 644614 355574 680058
rect 354954 644058 354986 644614
rect 355542 644058 355574 644614
rect 354954 608614 355574 644058
rect 354954 608058 354986 608614
rect 355542 608058 355574 608614
rect 354954 572614 355574 608058
rect 354954 572058 354986 572614
rect 355542 572058 355574 572614
rect 354954 536614 355574 572058
rect 354954 536058 354986 536614
rect 355542 536058 355574 536614
rect 354954 500614 355574 536058
rect 354954 500058 354986 500614
rect 355542 500058 355574 500614
rect 354954 500000 355574 500058
rect 361794 704838 362414 705830
rect 361794 704282 361826 704838
rect 362382 704282 362414 704838
rect 361794 687454 362414 704282
rect 361794 686898 361826 687454
rect 362382 686898 362414 687454
rect 361794 651454 362414 686898
rect 361794 650898 361826 651454
rect 362382 650898 362414 651454
rect 361794 615454 362414 650898
rect 361794 614898 361826 615454
rect 362382 614898 362414 615454
rect 361794 579454 362414 614898
rect 361794 578898 361826 579454
rect 362382 578898 362414 579454
rect 361794 543454 362414 578898
rect 361794 542898 361826 543454
rect 362382 542898 362414 543454
rect 361794 507454 362414 542898
rect 361794 506898 361826 507454
rect 362382 506898 362414 507454
rect 361794 500000 362414 506898
rect 365514 691174 366134 706202
rect 365514 690618 365546 691174
rect 366102 690618 366134 691174
rect 365514 655174 366134 690618
rect 365514 654618 365546 655174
rect 366102 654618 366134 655174
rect 365514 619174 366134 654618
rect 365514 618618 365546 619174
rect 366102 618618 366134 619174
rect 365514 583174 366134 618618
rect 365514 582618 365546 583174
rect 366102 582618 366134 583174
rect 365514 547174 366134 582618
rect 365514 546618 365546 547174
rect 366102 546618 366134 547174
rect 365514 511174 366134 546618
rect 365514 510618 365546 511174
rect 366102 510618 366134 511174
rect 365514 500000 366134 510618
rect 369234 694894 369854 708122
rect 369234 694338 369266 694894
rect 369822 694338 369854 694894
rect 369234 658894 369854 694338
rect 369234 658338 369266 658894
rect 369822 658338 369854 658894
rect 369234 622894 369854 658338
rect 369234 622338 369266 622894
rect 369822 622338 369854 622894
rect 369234 586894 369854 622338
rect 369234 586338 369266 586894
rect 369822 586338 369854 586894
rect 369234 550894 369854 586338
rect 369234 550338 369266 550894
rect 369822 550338 369854 550894
rect 369234 514894 369854 550338
rect 369234 514338 369266 514894
rect 369822 514338 369854 514894
rect 369234 500000 369854 514338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711002 390986 711558
rect 391542 711002 391574 711558
rect 387234 709638 387854 709670
rect 387234 709082 387266 709638
rect 387822 709082 387854 709638
rect 383514 707718 384134 707750
rect 383514 707162 383546 707718
rect 384102 707162 384134 707718
rect 372954 698058 372986 698614
rect 373542 698058 373574 698614
rect 372954 662614 373574 698058
rect 372954 662058 372986 662614
rect 373542 662058 373574 662614
rect 372954 626614 373574 662058
rect 372954 626058 372986 626614
rect 373542 626058 373574 626614
rect 372954 590614 373574 626058
rect 372954 590058 372986 590614
rect 373542 590058 373574 590614
rect 372954 554614 373574 590058
rect 372954 554058 372986 554614
rect 373542 554058 373574 554614
rect 372954 518614 373574 554058
rect 372954 518058 372986 518614
rect 373542 518058 373574 518614
rect 372954 500000 373574 518058
rect 379794 705798 380414 705830
rect 379794 705242 379826 705798
rect 380382 705242 380414 705798
rect 379794 669454 380414 705242
rect 379794 668898 379826 669454
rect 380382 668898 380414 669454
rect 379794 633454 380414 668898
rect 379794 632898 379826 633454
rect 380382 632898 380414 633454
rect 379794 597454 380414 632898
rect 379794 596898 379826 597454
rect 380382 596898 380414 597454
rect 379794 561454 380414 596898
rect 379794 560898 379826 561454
rect 380382 560898 380414 561454
rect 379794 525454 380414 560898
rect 379794 524898 379826 525454
rect 380382 524898 380414 525454
rect 379794 500000 380414 524898
rect 383514 673174 384134 707162
rect 383514 672618 383546 673174
rect 384102 672618 384134 673174
rect 383514 637174 384134 672618
rect 383514 636618 383546 637174
rect 384102 636618 384134 637174
rect 383514 601174 384134 636618
rect 383514 600618 383546 601174
rect 384102 600618 384134 601174
rect 383514 565174 384134 600618
rect 383514 564618 383546 565174
rect 384102 564618 384134 565174
rect 383514 529174 384134 564618
rect 383514 528618 383546 529174
rect 384102 528618 384134 529174
rect 383514 500000 384134 528618
rect 387234 676894 387854 709082
rect 387234 676338 387266 676894
rect 387822 676338 387854 676894
rect 387234 640894 387854 676338
rect 387234 640338 387266 640894
rect 387822 640338 387854 640894
rect 387234 604894 387854 640338
rect 387234 604338 387266 604894
rect 387822 604338 387854 604894
rect 387234 568894 387854 604338
rect 387234 568338 387266 568894
rect 387822 568338 387854 568894
rect 387234 532894 387854 568338
rect 387234 532338 387266 532894
rect 387822 532338 387854 532894
rect 387234 500000 387854 532338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710042 408986 710598
rect 409542 710042 409574 710598
rect 405234 708678 405854 709670
rect 405234 708122 405266 708678
rect 405822 708122 405854 708678
rect 401514 706758 402134 707750
rect 401514 706202 401546 706758
rect 402102 706202 402134 706758
rect 390954 680058 390986 680614
rect 391542 680058 391574 680614
rect 390954 644614 391574 680058
rect 390954 644058 390986 644614
rect 391542 644058 391574 644614
rect 390954 608614 391574 644058
rect 390954 608058 390986 608614
rect 391542 608058 391574 608614
rect 390954 572614 391574 608058
rect 390954 572058 390986 572614
rect 391542 572058 391574 572614
rect 390954 536614 391574 572058
rect 390954 536058 390986 536614
rect 391542 536058 391574 536614
rect 390954 500614 391574 536058
rect 390954 500058 390986 500614
rect 391542 500058 391574 500614
rect 390954 500000 391574 500058
rect 397794 704838 398414 705830
rect 397794 704282 397826 704838
rect 398382 704282 398414 704838
rect 397794 687454 398414 704282
rect 397794 686898 397826 687454
rect 398382 686898 398414 687454
rect 397794 651454 398414 686898
rect 397794 650898 397826 651454
rect 398382 650898 398414 651454
rect 397794 615454 398414 650898
rect 397794 614898 397826 615454
rect 398382 614898 398414 615454
rect 397794 579454 398414 614898
rect 397794 578898 397826 579454
rect 398382 578898 398414 579454
rect 397794 543454 398414 578898
rect 397794 542898 397826 543454
rect 398382 542898 398414 543454
rect 397794 507454 398414 542898
rect 397794 506898 397826 507454
rect 398382 506898 398414 507454
rect 397794 500000 398414 506898
rect 401514 691174 402134 706202
rect 401514 690618 401546 691174
rect 402102 690618 402134 691174
rect 401514 655174 402134 690618
rect 401514 654618 401546 655174
rect 402102 654618 402134 655174
rect 401514 619174 402134 654618
rect 401514 618618 401546 619174
rect 402102 618618 402134 619174
rect 401514 583174 402134 618618
rect 401514 582618 401546 583174
rect 402102 582618 402134 583174
rect 401514 547174 402134 582618
rect 401514 546618 401546 547174
rect 402102 546618 402134 547174
rect 401514 511174 402134 546618
rect 401514 510618 401546 511174
rect 402102 510618 402134 511174
rect 401514 500000 402134 510618
rect 405234 694894 405854 708122
rect 405234 694338 405266 694894
rect 405822 694338 405854 694894
rect 405234 658894 405854 694338
rect 405234 658338 405266 658894
rect 405822 658338 405854 658894
rect 405234 622894 405854 658338
rect 405234 622338 405266 622894
rect 405822 622338 405854 622894
rect 405234 586894 405854 622338
rect 405234 586338 405266 586894
rect 405822 586338 405854 586894
rect 405234 550894 405854 586338
rect 405234 550338 405266 550894
rect 405822 550338 405854 550894
rect 405234 514894 405854 550338
rect 405234 514338 405266 514894
rect 405822 514338 405854 514894
rect 405234 500000 405854 514338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711002 426986 711558
rect 427542 711002 427574 711558
rect 423234 709638 423854 709670
rect 423234 709082 423266 709638
rect 423822 709082 423854 709638
rect 419514 707718 420134 707750
rect 419514 707162 419546 707718
rect 420102 707162 420134 707718
rect 408954 698058 408986 698614
rect 409542 698058 409574 698614
rect 408954 662614 409574 698058
rect 408954 662058 408986 662614
rect 409542 662058 409574 662614
rect 408954 626614 409574 662058
rect 408954 626058 408986 626614
rect 409542 626058 409574 626614
rect 408954 590614 409574 626058
rect 408954 590058 408986 590614
rect 409542 590058 409574 590614
rect 408954 554614 409574 590058
rect 408954 554058 408986 554614
rect 409542 554058 409574 554614
rect 408954 518614 409574 554058
rect 408954 518058 408986 518614
rect 409542 518058 409574 518614
rect 408954 500000 409574 518058
rect 415794 705798 416414 705830
rect 415794 705242 415826 705798
rect 416382 705242 416414 705798
rect 415794 669454 416414 705242
rect 415794 668898 415826 669454
rect 416382 668898 416414 669454
rect 415794 633454 416414 668898
rect 415794 632898 415826 633454
rect 416382 632898 416414 633454
rect 415794 597454 416414 632898
rect 415794 596898 415826 597454
rect 416382 596898 416414 597454
rect 415794 561454 416414 596898
rect 415794 560898 415826 561454
rect 416382 560898 416414 561454
rect 415794 525454 416414 560898
rect 415794 524898 415826 525454
rect 416382 524898 416414 525454
rect 415794 500000 416414 524898
rect 419514 673174 420134 707162
rect 419514 672618 419546 673174
rect 420102 672618 420134 673174
rect 419514 637174 420134 672618
rect 419514 636618 419546 637174
rect 420102 636618 420134 637174
rect 419514 601174 420134 636618
rect 419514 600618 419546 601174
rect 420102 600618 420134 601174
rect 419514 565174 420134 600618
rect 419514 564618 419546 565174
rect 420102 564618 420134 565174
rect 419514 529174 420134 564618
rect 419514 528618 419546 529174
rect 420102 528618 420134 529174
rect 419514 500000 420134 528618
rect 423234 676894 423854 709082
rect 423234 676338 423266 676894
rect 423822 676338 423854 676894
rect 423234 640894 423854 676338
rect 423234 640338 423266 640894
rect 423822 640338 423854 640894
rect 423234 604894 423854 640338
rect 423234 604338 423266 604894
rect 423822 604338 423854 604894
rect 423234 568894 423854 604338
rect 423234 568338 423266 568894
rect 423822 568338 423854 568894
rect 423234 532894 423854 568338
rect 423234 532338 423266 532894
rect 423822 532338 423854 532894
rect 423234 500000 423854 532338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710042 444986 710598
rect 445542 710042 445574 710598
rect 441234 708678 441854 709670
rect 441234 708122 441266 708678
rect 441822 708122 441854 708678
rect 437514 706758 438134 707750
rect 437514 706202 437546 706758
rect 438102 706202 438134 706758
rect 426954 680058 426986 680614
rect 427542 680058 427574 680614
rect 426954 644614 427574 680058
rect 426954 644058 426986 644614
rect 427542 644058 427574 644614
rect 426954 608614 427574 644058
rect 426954 608058 426986 608614
rect 427542 608058 427574 608614
rect 426954 572614 427574 608058
rect 426954 572058 426986 572614
rect 427542 572058 427574 572614
rect 426954 536614 427574 572058
rect 426954 536058 426986 536614
rect 427542 536058 427574 536614
rect 426954 500614 427574 536058
rect 426954 500058 426986 500614
rect 427542 500058 427574 500614
rect 426954 500000 427574 500058
rect 433794 704838 434414 705830
rect 433794 704282 433826 704838
rect 434382 704282 434414 704838
rect 433794 687454 434414 704282
rect 433794 686898 433826 687454
rect 434382 686898 434414 687454
rect 433794 651454 434414 686898
rect 433794 650898 433826 651454
rect 434382 650898 434414 651454
rect 433794 615454 434414 650898
rect 433794 614898 433826 615454
rect 434382 614898 434414 615454
rect 433794 579454 434414 614898
rect 433794 578898 433826 579454
rect 434382 578898 434414 579454
rect 433794 543454 434414 578898
rect 433794 542898 433826 543454
rect 434382 542898 434414 543454
rect 433794 507454 434414 542898
rect 433794 506898 433826 507454
rect 434382 506898 434414 507454
rect 433794 500000 434414 506898
rect 437514 691174 438134 706202
rect 437514 690618 437546 691174
rect 438102 690618 438134 691174
rect 437514 655174 438134 690618
rect 437514 654618 437546 655174
rect 438102 654618 438134 655174
rect 437514 619174 438134 654618
rect 437514 618618 437546 619174
rect 438102 618618 438134 619174
rect 437514 583174 438134 618618
rect 437514 582618 437546 583174
rect 438102 582618 438134 583174
rect 437514 547174 438134 582618
rect 437514 546618 437546 547174
rect 438102 546618 438134 547174
rect 437514 511174 438134 546618
rect 437514 510618 437546 511174
rect 438102 510618 438134 511174
rect 400443 497588 400509 497589
rect 400443 497524 400444 497588
rect 400508 497524 400509 497588
rect 400443 497523 400509 497524
rect 418107 497588 418173 497589
rect 418107 497524 418108 497588
rect 418172 497524 418173 497588
rect 418107 497523 418173 497524
rect 238523 497452 238589 497453
rect 238523 497388 238524 497452
rect 238588 497388 238589 497452
rect 238523 497387 238589 497388
rect 254899 497452 254965 497453
rect 254899 497388 254900 497452
rect 254964 497388 254965 497452
rect 254899 497387 254965 497388
rect 262075 497452 262141 497453
rect 262075 497388 262076 497452
rect 262140 497388 262141 497452
rect 265019 497452 265085 497453
rect 265019 497450 265020 497452
rect 262075 497387 262141 497388
rect 264654 497390 265020 497450
rect 236683 318884 236749 318885
rect 236683 318820 236684 318884
rect 236748 318820 236749 318884
rect 236683 318819 236749 318820
rect 236499 266388 236565 266389
rect 236499 266324 236500 266388
rect 236564 266324 236565 266388
rect 236499 266323 236565 266324
rect 235794 236898 235826 237454
rect 236382 236898 236414 237454
rect 235794 201454 236414 236898
rect 235794 200898 235826 201454
rect 236382 200898 236414 201454
rect 235794 165454 236414 200898
rect 235794 164898 235826 165454
rect 236382 164898 236414 165454
rect 235794 129454 236414 164898
rect 235794 128898 235826 129454
rect 236382 128898 236414 129454
rect 235794 93454 236414 128898
rect 235794 92898 235826 93454
rect 236382 92898 236414 93454
rect 233739 84284 233805 84285
rect 233739 84220 233740 84284
rect 233804 84220 233805 84284
rect 233739 84219 233805 84220
rect 228954 50058 228986 50614
rect 229542 50058 229574 50614
rect 228954 14614 229574 50058
rect 228954 14058 228986 14614
rect 229542 14058 229574 14614
rect 210954 -7622 210986 -7066
rect 211542 -7622 211574 -7066
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 92898
rect 235794 56898 235826 57454
rect 236382 56898 236414 57454
rect 235794 21454 236414 56898
rect 238526 31925 238586 497387
rect 254902 496909 254962 497387
rect 262078 497045 262138 497387
rect 264654 497317 264714 497390
rect 265019 497388 265020 497390
rect 265084 497388 265085 497452
rect 265019 497387 265085 497388
rect 264651 497316 264717 497317
rect 264651 497252 264652 497316
rect 264716 497252 264717 497316
rect 264651 497251 264717 497252
rect 262075 497044 262141 497045
rect 262075 496980 262076 497044
rect 262140 496980 262141 497044
rect 262075 496979 262141 496980
rect 254899 496908 254965 496909
rect 254899 496844 254900 496908
rect 254964 496844 254965 496908
rect 254899 496843 254965 496844
rect 400446 496229 400506 497523
rect 400443 496228 400509 496229
rect 400443 496164 400444 496228
rect 400508 496164 400509 496228
rect 400443 496163 400509 496164
rect 418110 496093 418170 497523
rect 423995 497452 424061 497453
rect 423995 497388 423996 497452
rect 424060 497388 424061 497452
rect 423995 497387 424061 497388
rect 425099 497452 425165 497453
rect 425099 497388 425100 497452
rect 425164 497388 425165 497452
rect 425099 497387 425165 497388
rect 426387 497452 426453 497453
rect 426387 497388 426388 497452
rect 426452 497388 426453 497452
rect 426387 497387 426453 497388
rect 427859 497452 427925 497453
rect 427859 497388 427860 497452
rect 427924 497388 427925 497452
rect 427859 497387 427925 497388
rect 429147 497452 429213 497453
rect 429147 497388 429148 497452
rect 429212 497388 429213 497452
rect 429147 497387 429213 497388
rect 433379 497452 433445 497453
rect 433379 497388 433380 497452
rect 433444 497388 433445 497452
rect 433379 497387 433445 497388
rect 418107 496092 418173 496093
rect 418107 496028 418108 496092
rect 418172 496028 418173 496092
rect 418107 496027 418173 496028
rect 254568 489454 254888 489486
rect 254568 489218 254610 489454
rect 254846 489218 254888 489454
rect 254568 489134 254888 489218
rect 254568 488898 254610 489134
rect 254846 488898 254888 489134
rect 254568 488866 254888 488898
rect 285288 489454 285608 489486
rect 285288 489218 285330 489454
rect 285566 489218 285608 489454
rect 285288 489134 285608 489218
rect 285288 488898 285330 489134
rect 285566 488898 285608 489134
rect 285288 488866 285608 488898
rect 316008 489454 316328 489486
rect 316008 489218 316050 489454
rect 316286 489218 316328 489454
rect 316008 489134 316328 489218
rect 316008 488898 316050 489134
rect 316286 488898 316328 489134
rect 316008 488866 316328 488898
rect 346728 489454 347048 489486
rect 346728 489218 346770 489454
rect 347006 489218 347048 489454
rect 346728 489134 347048 489218
rect 346728 488898 346770 489134
rect 347006 488898 347048 489134
rect 346728 488866 347048 488898
rect 377448 489454 377768 489486
rect 377448 489218 377490 489454
rect 377726 489218 377768 489454
rect 377448 489134 377768 489218
rect 377448 488898 377490 489134
rect 377726 488898 377768 489134
rect 377448 488866 377768 488898
rect 408168 489454 408488 489486
rect 408168 489218 408210 489454
rect 408446 489218 408488 489454
rect 408168 489134 408488 489218
rect 408168 488898 408210 489134
rect 408446 488898 408488 489134
rect 408168 488866 408488 488898
rect 239208 471454 239528 471486
rect 239208 471218 239250 471454
rect 239486 471218 239528 471454
rect 239208 471134 239528 471218
rect 239208 470898 239250 471134
rect 239486 470898 239528 471134
rect 239208 470866 239528 470898
rect 269928 471454 270248 471486
rect 269928 471218 269970 471454
rect 270206 471218 270248 471454
rect 269928 471134 270248 471218
rect 269928 470898 269970 471134
rect 270206 470898 270248 471134
rect 269928 470866 270248 470898
rect 300648 471454 300968 471486
rect 300648 471218 300690 471454
rect 300926 471218 300968 471454
rect 300648 471134 300968 471218
rect 300648 470898 300690 471134
rect 300926 470898 300968 471134
rect 300648 470866 300968 470898
rect 331368 471454 331688 471486
rect 331368 471218 331410 471454
rect 331646 471218 331688 471454
rect 331368 471134 331688 471218
rect 331368 470898 331410 471134
rect 331646 470898 331688 471134
rect 331368 470866 331688 470898
rect 362088 471454 362408 471486
rect 362088 471218 362130 471454
rect 362366 471218 362408 471454
rect 362088 471134 362408 471218
rect 362088 470898 362130 471134
rect 362366 470898 362408 471134
rect 362088 470866 362408 470898
rect 392808 471454 393128 471486
rect 392808 471218 392850 471454
rect 393086 471218 393128 471454
rect 392808 471134 393128 471218
rect 392808 470898 392850 471134
rect 393086 470898 393128 471134
rect 392808 470866 393128 470898
rect 423528 471454 423848 471486
rect 423528 471218 423570 471454
rect 423806 471218 423848 471454
rect 423528 471134 423848 471218
rect 423528 470898 423570 471134
rect 423806 470898 423848 471134
rect 423528 470866 423848 470898
rect 254568 453454 254888 453486
rect 254568 453218 254610 453454
rect 254846 453218 254888 453454
rect 254568 453134 254888 453218
rect 254568 452898 254610 453134
rect 254846 452898 254888 453134
rect 254568 452866 254888 452898
rect 285288 453454 285608 453486
rect 285288 453218 285330 453454
rect 285566 453218 285608 453454
rect 285288 453134 285608 453218
rect 285288 452898 285330 453134
rect 285566 452898 285608 453134
rect 285288 452866 285608 452898
rect 316008 453454 316328 453486
rect 316008 453218 316050 453454
rect 316286 453218 316328 453454
rect 316008 453134 316328 453218
rect 316008 452898 316050 453134
rect 316286 452898 316328 453134
rect 316008 452866 316328 452898
rect 346728 453454 347048 453486
rect 346728 453218 346770 453454
rect 347006 453218 347048 453454
rect 346728 453134 347048 453218
rect 346728 452898 346770 453134
rect 347006 452898 347048 453134
rect 346728 452866 347048 452898
rect 377448 453454 377768 453486
rect 377448 453218 377490 453454
rect 377726 453218 377768 453454
rect 377448 453134 377768 453218
rect 377448 452898 377490 453134
rect 377726 452898 377768 453134
rect 377448 452866 377768 452898
rect 408168 453454 408488 453486
rect 408168 453218 408210 453454
rect 408446 453218 408488 453454
rect 408168 453134 408488 453218
rect 408168 452898 408210 453134
rect 408446 452898 408488 453134
rect 408168 452866 408488 452898
rect 239208 435454 239528 435486
rect 239208 435218 239250 435454
rect 239486 435218 239528 435454
rect 239208 435134 239528 435218
rect 239208 434898 239250 435134
rect 239486 434898 239528 435134
rect 239208 434866 239528 434898
rect 269928 435454 270248 435486
rect 269928 435218 269970 435454
rect 270206 435218 270248 435454
rect 269928 435134 270248 435218
rect 269928 434898 269970 435134
rect 270206 434898 270248 435134
rect 269928 434866 270248 434898
rect 300648 435454 300968 435486
rect 300648 435218 300690 435454
rect 300926 435218 300968 435454
rect 300648 435134 300968 435218
rect 300648 434898 300690 435134
rect 300926 434898 300968 435134
rect 300648 434866 300968 434898
rect 331368 435454 331688 435486
rect 331368 435218 331410 435454
rect 331646 435218 331688 435454
rect 331368 435134 331688 435218
rect 331368 434898 331410 435134
rect 331646 434898 331688 435134
rect 331368 434866 331688 434898
rect 362088 435454 362408 435486
rect 362088 435218 362130 435454
rect 362366 435218 362408 435454
rect 362088 435134 362408 435218
rect 362088 434898 362130 435134
rect 362366 434898 362408 435134
rect 362088 434866 362408 434898
rect 392808 435454 393128 435486
rect 392808 435218 392850 435454
rect 393086 435218 393128 435454
rect 392808 435134 393128 435218
rect 392808 434898 392850 435134
rect 393086 434898 393128 435134
rect 392808 434866 393128 434898
rect 423528 435454 423848 435486
rect 423528 435218 423570 435454
rect 423806 435218 423848 435454
rect 423528 435134 423848 435218
rect 423528 434898 423570 435134
rect 423806 434898 423848 435134
rect 423528 434866 423848 434898
rect 254568 417454 254888 417486
rect 254568 417218 254610 417454
rect 254846 417218 254888 417454
rect 254568 417134 254888 417218
rect 254568 416898 254610 417134
rect 254846 416898 254888 417134
rect 254568 416866 254888 416898
rect 285288 417454 285608 417486
rect 285288 417218 285330 417454
rect 285566 417218 285608 417454
rect 285288 417134 285608 417218
rect 285288 416898 285330 417134
rect 285566 416898 285608 417134
rect 285288 416866 285608 416898
rect 316008 417454 316328 417486
rect 316008 417218 316050 417454
rect 316286 417218 316328 417454
rect 316008 417134 316328 417218
rect 316008 416898 316050 417134
rect 316286 416898 316328 417134
rect 316008 416866 316328 416898
rect 346728 417454 347048 417486
rect 346728 417218 346770 417454
rect 347006 417218 347048 417454
rect 346728 417134 347048 417218
rect 346728 416898 346770 417134
rect 347006 416898 347048 417134
rect 346728 416866 347048 416898
rect 377448 417454 377768 417486
rect 377448 417218 377490 417454
rect 377726 417218 377768 417454
rect 377448 417134 377768 417218
rect 377448 416898 377490 417134
rect 377726 416898 377768 417134
rect 377448 416866 377768 416898
rect 408168 417454 408488 417486
rect 408168 417218 408210 417454
rect 408446 417218 408488 417454
rect 408168 417134 408488 417218
rect 408168 416898 408210 417134
rect 408446 416898 408488 417134
rect 408168 416866 408488 416898
rect 239208 399454 239528 399486
rect 239208 399218 239250 399454
rect 239486 399218 239528 399454
rect 239208 399134 239528 399218
rect 239208 398898 239250 399134
rect 239486 398898 239528 399134
rect 239208 398866 239528 398898
rect 269928 399454 270248 399486
rect 269928 399218 269970 399454
rect 270206 399218 270248 399454
rect 269928 399134 270248 399218
rect 269928 398898 269970 399134
rect 270206 398898 270248 399134
rect 269928 398866 270248 398898
rect 300648 399454 300968 399486
rect 300648 399218 300690 399454
rect 300926 399218 300968 399454
rect 300648 399134 300968 399218
rect 300648 398898 300690 399134
rect 300926 398898 300968 399134
rect 300648 398866 300968 398898
rect 331368 399454 331688 399486
rect 331368 399218 331410 399454
rect 331646 399218 331688 399454
rect 331368 399134 331688 399218
rect 331368 398898 331410 399134
rect 331646 398898 331688 399134
rect 331368 398866 331688 398898
rect 362088 399454 362408 399486
rect 362088 399218 362130 399454
rect 362366 399218 362408 399454
rect 362088 399134 362408 399218
rect 362088 398898 362130 399134
rect 362366 398898 362408 399134
rect 362088 398866 362408 398898
rect 392808 399454 393128 399486
rect 392808 399218 392850 399454
rect 393086 399218 393128 399454
rect 392808 399134 393128 399218
rect 392808 398898 392850 399134
rect 393086 398898 393128 399134
rect 392808 398866 393128 398898
rect 423528 399454 423848 399486
rect 423528 399218 423570 399454
rect 423806 399218 423848 399454
rect 423528 399134 423848 399218
rect 423528 398898 423570 399134
rect 423806 398898 423848 399134
rect 423528 398866 423848 398898
rect 254568 381454 254888 381486
rect 254568 381218 254610 381454
rect 254846 381218 254888 381454
rect 254568 381134 254888 381218
rect 254568 380898 254610 381134
rect 254846 380898 254888 381134
rect 254568 380866 254888 380898
rect 285288 381454 285608 381486
rect 285288 381218 285330 381454
rect 285566 381218 285608 381454
rect 285288 381134 285608 381218
rect 285288 380898 285330 381134
rect 285566 380898 285608 381134
rect 285288 380866 285608 380898
rect 316008 381454 316328 381486
rect 316008 381218 316050 381454
rect 316286 381218 316328 381454
rect 316008 381134 316328 381218
rect 316008 380898 316050 381134
rect 316286 380898 316328 381134
rect 316008 380866 316328 380898
rect 346728 381454 347048 381486
rect 346728 381218 346770 381454
rect 347006 381218 347048 381454
rect 346728 381134 347048 381218
rect 346728 380898 346770 381134
rect 347006 380898 347048 381134
rect 346728 380866 347048 380898
rect 377448 381454 377768 381486
rect 377448 381218 377490 381454
rect 377726 381218 377768 381454
rect 377448 381134 377768 381218
rect 377448 380898 377490 381134
rect 377726 380898 377768 381134
rect 377448 380866 377768 380898
rect 408168 381454 408488 381486
rect 408168 381218 408210 381454
rect 408446 381218 408488 381454
rect 408168 381134 408488 381218
rect 408168 380898 408210 381134
rect 408446 380898 408488 381134
rect 408168 380866 408488 380898
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 300648 363454 300968 363486
rect 300648 363218 300690 363454
rect 300926 363218 300968 363454
rect 300648 363134 300968 363218
rect 300648 362898 300690 363134
rect 300926 362898 300968 363134
rect 300648 362866 300968 362898
rect 331368 363454 331688 363486
rect 331368 363218 331410 363454
rect 331646 363218 331688 363454
rect 331368 363134 331688 363218
rect 331368 362898 331410 363134
rect 331646 362898 331688 363134
rect 331368 362866 331688 362898
rect 362088 363454 362408 363486
rect 362088 363218 362130 363454
rect 362366 363218 362408 363454
rect 362088 363134 362408 363218
rect 362088 362898 362130 363134
rect 362366 362898 362408 363134
rect 362088 362866 362408 362898
rect 392808 363454 393128 363486
rect 392808 363218 392850 363454
rect 393086 363218 393128 363454
rect 392808 363134 393128 363218
rect 392808 362898 392850 363134
rect 393086 362898 393128 363134
rect 392808 362866 393128 362898
rect 423528 363454 423848 363486
rect 423528 363218 423570 363454
rect 423806 363218 423848 363454
rect 423528 363134 423848 363218
rect 423528 362898 423570 363134
rect 423806 362898 423848 363134
rect 423528 362866 423848 362898
rect 254568 345454 254888 345486
rect 254568 345218 254610 345454
rect 254846 345218 254888 345454
rect 254568 345134 254888 345218
rect 254568 344898 254610 345134
rect 254846 344898 254888 345134
rect 254568 344866 254888 344898
rect 285288 345454 285608 345486
rect 285288 345218 285330 345454
rect 285566 345218 285608 345454
rect 285288 345134 285608 345218
rect 285288 344898 285330 345134
rect 285566 344898 285608 345134
rect 285288 344866 285608 344898
rect 316008 345454 316328 345486
rect 316008 345218 316050 345454
rect 316286 345218 316328 345454
rect 316008 345134 316328 345218
rect 316008 344898 316050 345134
rect 316286 344898 316328 345134
rect 316008 344866 316328 344898
rect 346728 345454 347048 345486
rect 346728 345218 346770 345454
rect 347006 345218 347048 345454
rect 346728 345134 347048 345218
rect 346728 344898 346770 345134
rect 347006 344898 347048 345134
rect 346728 344866 347048 344898
rect 377448 345454 377768 345486
rect 377448 345218 377490 345454
rect 377726 345218 377768 345454
rect 377448 345134 377768 345218
rect 377448 344898 377490 345134
rect 377726 344898 377768 345134
rect 377448 344866 377768 344898
rect 408168 345454 408488 345486
rect 408168 345218 408210 345454
rect 408446 345218 408488 345454
rect 408168 345134 408488 345218
rect 408168 344898 408210 345134
rect 408446 344898 408488 345134
rect 408168 344866 408488 344898
rect 239514 313174 240134 336000
rect 239514 312618 239546 313174
rect 240102 312618 240134 313174
rect 239514 277174 240134 312618
rect 239514 276618 239546 277174
rect 240102 276618 240134 277174
rect 239514 241174 240134 276618
rect 239514 240618 239546 241174
rect 240102 240618 240134 241174
rect 239514 205174 240134 240618
rect 239514 204618 239546 205174
rect 240102 204618 240134 205174
rect 239514 169174 240134 204618
rect 239514 168618 239546 169174
rect 240102 168618 240134 169174
rect 239514 133174 240134 168618
rect 239514 132618 239546 133174
rect 240102 132618 240134 133174
rect 239514 97174 240134 132618
rect 239514 96618 239546 97174
rect 240102 96618 240134 97174
rect 239514 61174 240134 96618
rect 239514 60618 239546 61174
rect 240102 60618 240134 61174
rect 238523 31924 238589 31925
rect 238523 31860 238524 31924
rect 238588 31860 238589 31924
rect 238523 31859 238589 31860
rect 235794 20898 235826 21454
rect 236382 20898 236414 21454
rect 235794 -1306 236414 20898
rect 235794 -1862 235826 -1306
rect 236382 -1862 236414 -1306
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 60618
rect 239514 24618 239546 25174
rect 240102 24618 240134 25174
rect 239514 -3226 240134 24618
rect 239514 -3782 239546 -3226
rect 240102 -3782 240134 -3226
rect 239514 -3814 240134 -3782
rect 243234 316894 243854 336000
rect 243234 316338 243266 316894
rect 243822 316338 243854 316894
rect 243234 280894 243854 316338
rect 243234 280338 243266 280894
rect 243822 280338 243854 280894
rect 243234 244894 243854 280338
rect 243234 244338 243266 244894
rect 243822 244338 243854 244894
rect 243234 208894 243854 244338
rect 243234 208338 243266 208894
rect 243822 208338 243854 208894
rect 243234 172894 243854 208338
rect 243234 172338 243266 172894
rect 243822 172338 243854 172894
rect 243234 136894 243854 172338
rect 243234 136338 243266 136894
rect 243822 136338 243854 136894
rect 243234 100894 243854 136338
rect 243234 100338 243266 100894
rect 243822 100338 243854 100894
rect 243234 64894 243854 100338
rect 243234 64338 243266 64894
rect 243822 64338 243854 64894
rect 243234 28894 243854 64338
rect 243234 28338 243266 28894
rect 243822 28338 243854 28894
rect 243234 -5146 243854 28338
rect 243234 -5702 243266 -5146
rect 243822 -5702 243854 -5146
rect 243234 -5734 243854 -5702
rect 246954 320614 247574 336000
rect 246954 320058 246986 320614
rect 247542 320058 247574 320614
rect 246954 284614 247574 320058
rect 246954 284058 246986 284614
rect 247542 284058 247574 284614
rect 246954 248614 247574 284058
rect 246954 248058 246986 248614
rect 247542 248058 247574 248614
rect 246954 212614 247574 248058
rect 246954 212058 246986 212614
rect 247542 212058 247574 212614
rect 246954 176614 247574 212058
rect 246954 176058 246986 176614
rect 247542 176058 247574 176614
rect 246954 140614 247574 176058
rect 246954 140058 246986 140614
rect 247542 140058 247574 140614
rect 246954 104614 247574 140058
rect 246954 104058 246986 104614
rect 247542 104058 247574 104614
rect 246954 68614 247574 104058
rect 246954 68058 246986 68614
rect 247542 68058 247574 68614
rect 246954 32614 247574 68058
rect 246954 32058 246986 32614
rect 247542 32058 247574 32614
rect 228954 -6662 228986 -6106
rect 229542 -6662 229574 -6106
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 327454 254414 336000
rect 253794 326898 253826 327454
rect 254382 326898 254414 327454
rect 253794 291454 254414 326898
rect 253794 290898 253826 291454
rect 254382 290898 254414 291454
rect 253794 255454 254414 290898
rect 253794 254898 253826 255454
rect 254382 254898 254414 255454
rect 253794 219454 254414 254898
rect 253794 218898 253826 219454
rect 254382 218898 254414 219454
rect 253794 183454 254414 218898
rect 253794 182898 253826 183454
rect 254382 182898 254414 183454
rect 253794 147454 254414 182898
rect 253794 146898 253826 147454
rect 254382 146898 254414 147454
rect 253794 111454 254414 146898
rect 253794 110898 253826 111454
rect 254382 110898 254414 111454
rect 253794 75454 254414 110898
rect 253794 74898 253826 75454
rect 254382 74898 254414 75454
rect 253794 39454 254414 74898
rect 253794 38898 253826 39454
rect 254382 38898 254414 39454
rect 253794 3454 254414 38898
rect 253794 2898 253826 3454
rect 254382 2898 254414 3454
rect 253794 -346 254414 2898
rect 253794 -902 253826 -346
rect 254382 -902 254414 -346
rect 253794 -1894 254414 -902
rect 257514 331174 258134 336000
rect 257514 330618 257546 331174
rect 258102 330618 258134 331174
rect 257514 295174 258134 330618
rect 257514 294618 257546 295174
rect 258102 294618 258134 295174
rect 257514 259174 258134 294618
rect 257514 258618 257546 259174
rect 258102 258618 258134 259174
rect 257514 223174 258134 258618
rect 257514 222618 257546 223174
rect 258102 222618 258134 223174
rect 257514 187174 258134 222618
rect 257514 186618 257546 187174
rect 258102 186618 258134 187174
rect 257514 151174 258134 186618
rect 257514 150618 257546 151174
rect 258102 150618 258134 151174
rect 257514 115174 258134 150618
rect 257514 114618 257546 115174
rect 258102 114618 258134 115174
rect 257514 79174 258134 114618
rect 257514 78618 257546 79174
rect 258102 78618 258134 79174
rect 257514 43174 258134 78618
rect 257514 42618 257546 43174
rect 258102 42618 258134 43174
rect 257514 7174 258134 42618
rect 257514 6618 257546 7174
rect 258102 6618 258134 7174
rect 257514 -2266 258134 6618
rect 257514 -2822 257546 -2266
rect 258102 -2822 258134 -2266
rect 257514 -3814 258134 -2822
rect 261234 334894 261854 336000
rect 261234 334338 261266 334894
rect 261822 334338 261854 334894
rect 261234 298894 261854 334338
rect 261234 298338 261266 298894
rect 261822 298338 261854 298894
rect 261234 262894 261854 298338
rect 261234 262338 261266 262894
rect 261822 262338 261854 262894
rect 261234 226894 261854 262338
rect 261234 226338 261266 226894
rect 261822 226338 261854 226894
rect 261234 190894 261854 226338
rect 261234 190338 261266 190894
rect 261822 190338 261854 190894
rect 261234 154894 261854 190338
rect 261234 154338 261266 154894
rect 261822 154338 261854 154894
rect 261234 118894 261854 154338
rect 261234 118338 261266 118894
rect 261822 118338 261854 118894
rect 261234 82894 261854 118338
rect 261234 82338 261266 82894
rect 261822 82338 261854 82894
rect 261234 46894 261854 82338
rect 261234 46338 261266 46894
rect 261822 46338 261854 46894
rect 261234 10894 261854 46338
rect 261234 10338 261266 10894
rect 261822 10338 261854 10894
rect 261234 -4186 261854 10338
rect 261234 -4742 261266 -4186
rect 261822 -4742 261854 -4186
rect 261234 -5734 261854 -4742
rect 264954 302614 265574 336000
rect 264954 302058 264986 302614
rect 265542 302058 265574 302614
rect 264954 266614 265574 302058
rect 264954 266058 264986 266614
rect 265542 266058 265574 266614
rect 264954 230614 265574 266058
rect 264954 230058 264986 230614
rect 265542 230058 265574 230614
rect 264954 194614 265574 230058
rect 264954 194058 264986 194614
rect 265542 194058 265574 194614
rect 264954 158614 265574 194058
rect 264954 158058 264986 158614
rect 265542 158058 265574 158614
rect 264954 122614 265574 158058
rect 264954 122058 264986 122614
rect 265542 122058 265574 122614
rect 264954 86614 265574 122058
rect 264954 86058 264986 86614
rect 265542 86058 265574 86614
rect 264954 50614 265574 86058
rect 264954 50058 264986 50614
rect 265542 50058 265574 50614
rect 264954 14614 265574 50058
rect 264954 14058 264986 14614
rect 265542 14058 265574 14614
rect 246954 -7622 246986 -7066
rect 247542 -7622 247574 -7066
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 309454 272414 336000
rect 271794 308898 271826 309454
rect 272382 308898 272414 309454
rect 271794 273454 272414 308898
rect 271794 272898 271826 273454
rect 272382 272898 272414 273454
rect 271794 237454 272414 272898
rect 271794 236898 271826 237454
rect 272382 236898 272414 237454
rect 271794 201454 272414 236898
rect 271794 200898 271826 201454
rect 272382 200898 272414 201454
rect 271794 165454 272414 200898
rect 271794 164898 271826 165454
rect 272382 164898 272414 165454
rect 271794 129454 272414 164898
rect 271794 128898 271826 129454
rect 272382 128898 272414 129454
rect 271794 93454 272414 128898
rect 271794 92898 271826 93454
rect 272382 92898 272414 93454
rect 271794 57454 272414 92898
rect 271794 56898 271826 57454
rect 272382 56898 272414 57454
rect 271794 21454 272414 56898
rect 271794 20898 271826 21454
rect 272382 20898 272414 21454
rect 271794 -1306 272414 20898
rect 271794 -1862 271826 -1306
rect 272382 -1862 272414 -1306
rect 271794 -1894 272414 -1862
rect 275514 313174 276134 336000
rect 275514 312618 275546 313174
rect 276102 312618 276134 313174
rect 275514 277174 276134 312618
rect 275514 276618 275546 277174
rect 276102 276618 276134 277174
rect 275514 241174 276134 276618
rect 275514 240618 275546 241174
rect 276102 240618 276134 241174
rect 275514 205174 276134 240618
rect 275514 204618 275546 205174
rect 276102 204618 276134 205174
rect 275514 169174 276134 204618
rect 275514 168618 275546 169174
rect 276102 168618 276134 169174
rect 275514 133174 276134 168618
rect 275514 132618 275546 133174
rect 276102 132618 276134 133174
rect 275514 97174 276134 132618
rect 275514 96618 275546 97174
rect 276102 96618 276134 97174
rect 275514 61174 276134 96618
rect 275514 60618 275546 61174
rect 276102 60618 276134 61174
rect 275514 25174 276134 60618
rect 275514 24618 275546 25174
rect 276102 24618 276134 25174
rect 275514 -3226 276134 24618
rect 275514 -3782 275546 -3226
rect 276102 -3782 276134 -3226
rect 275514 -3814 276134 -3782
rect 279234 316894 279854 336000
rect 279234 316338 279266 316894
rect 279822 316338 279854 316894
rect 279234 280894 279854 316338
rect 279234 280338 279266 280894
rect 279822 280338 279854 280894
rect 279234 244894 279854 280338
rect 279234 244338 279266 244894
rect 279822 244338 279854 244894
rect 279234 208894 279854 244338
rect 279234 208338 279266 208894
rect 279822 208338 279854 208894
rect 279234 172894 279854 208338
rect 279234 172338 279266 172894
rect 279822 172338 279854 172894
rect 279234 136894 279854 172338
rect 279234 136338 279266 136894
rect 279822 136338 279854 136894
rect 279234 100894 279854 136338
rect 279234 100338 279266 100894
rect 279822 100338 279854 100894
rect 279234 64894 279854 100338
rect 279234 64338 279266 64894
rect 279822 64338 279854 64894
rect 279234 28894 279854 64338
rect 279234 28338 279266 28894
rect 279822 28338 279854 28894
rect 279234 -5146 279854 28338
rect 279234 -5702 279266 -5146
rect 279822 -5702 279854 -5146
rect 279234 -5734 279854 -5702
rect 282954 320614 283574 336000
rect 282954 320058 282986 320614
rect 283542 320058 283574 320614
rect 282954 284614 283574 320058
rect 282954 284058 282986 284614
rect 283542 284058 283574 284614
rect 282954 248614 283574 284058
rect 282954 248058 282986 248614
rect 283542 248058 283574 248614
rect 282954 212614 283574 248058
rect 282954 212058 282986 212614
rect 283542 212058 283574 212614
rect 282954 176614 283574 212058
rect 282954 176058 282986 176614
rect 283542 176058 283574 176614
rect 282954 140614 283574 176058
rect 282954 140058 282986 140614
rect 283542 140058 283574 140614
rect 282954 104614 283574 140058
rect 282954 104058 282986 104614
rect 283542 104058 283574 104614
rect 282954 68614 283574 104058
rect 282954 68058 282986 68614
rect 283542 68058 283574 68614
rect 282954 32614 283574 68058
rect 282954 32058 282986 32614
rect 283542 32058 283574 32614
rect 264954 -6662 264986 -6106
rect 265542 -6662 265574 -6106
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 327454 290414 336000
rect 289794 326898 289826 327454
rect 290382 326898 290414 327454
rect 289794 291454 290414 326898
rect 289794 290898 289826 291454
rect 290382 290898 290414 291454
rect 289794 255454 290414 290898
rect 289794 254898 289826 255454
rect 290382 254898 290414 255454
rect 289794 219454 290414 254898
rect 289794 218898 289826 219454
rect 290382 218898 290414 219454
rect 289794 183454 290414 218898
rect 289794 182898 289826 183454
rect 290382 182898 290414 183454
rect 289794 147454 290414 182898
rect 289794 146898 289826 147454
rect 290382 146898 290414 147454
rect 289794 111454 290414 146898
rect 289794 110898 289826 111454
rect 290382 110898 290414 111454
rect 289794 75454 290414 110898
rect 289794 74898 289826 75454
rect 290382 74898 290414 75454
rect 289794 39454 290414 74898
rect 289794 38898 289826 39454
rect 290382 38898 290414 39454
rect 289794 3454 290414 38898
rect 289794 2898 289826 3454
rect 290382 2898 290414 3454
rect 289794 -346 290414 2898
rect 289794 -902 289826 -346
rect 290382 -902 290414 -346
rect 289794 -1894 290414 -902
rect 293514 331174 294134 336000
rect 293514 330618 293546 331174
rect 294102 330618 294134 331174
rect 293514 295174 294134 330618
rect 293514 294618 293546 295174
rect 294102 294618 294134 295174
rect 293514 259174 294134 294618
rect 293514 258618 293546 259174
rect 294102 258618 294134 259174
rect 293514 223174 294134 258618
rect 293514 222618 293546 223174
rect 294102 222618 294134 223174
rect 293514 187174 294134 222618
rect 293514 186618 293546 187174
rect 294102 186618 294134 187174
rect 293514 151174 294134 186618
rect 293514 150618 293546 151174
rect 294102 150618 294134 151174
rect 293514 115174 294134 150618
rect 293514 114618 293546 115174
rect 294102 114618 294134 115174
rect 293514 79174 294134 114618
rect 293514 78618 293546 79174
rect 294102 78618 294134 79174
rect 293514 43174 294134 78618
rect 293514 42618 293546 43174
rect 294102 42618 294134 43174
rect 293514 7174 294134 42618
rect 293514 6618 293546 7174
rect 294102 6618 294134 7174
rect 293514 -2266 294134 6618
rect 293514 -2822 293546 -2266
rect 294102 -2822 294134 -2266
rect 293514 -3814 294134 -2822
rect 297234 334894 297854 336000
rect 297234 334338 297266 334894
rect 297822 334338 297854 334894
rect 297234 298894 297854 334338
rect 297234 298338 297266 298894
rect 297822 298338 297854 298894
rect 297234 262894 297854 298338
rect 297234 262338 297266 262894
rect 297822 262338 297854 262894
rect 297234 226894 297854 262338
rect 297234 226338 297266 226894
rect 297822 226338 297854 226894
rect 297234 190894 297854 226338
rect 297234 190338 297266 190894
rect 297822 190338 297854 190894
rect 297234 154894 297854 190338
rect 297234 154338 297266 154894
rect 297822 154338 297854 154894
rect 297234 118894 297854 154338
rect 297234 118338 297266 118894
rect 297822 118338 297854 118894
rect 297234 82894 297854 118338
rect 297234 82338 297266 82894
rect 297822 82338 297854 82894
rect 297234 46894 297854 82338
rect 297234 46338 297266 46894
rect 297822 46338 297854 46894
rect 297234 10894 297854 46338
rect 297234 10338 297266 10894
rect 297822 10338 297854 10894
rect 297234 -4186 297854 10338
rect 297234 -4742 297266 -4186
rect 297822 -4742 297854 -4186
rect 297234 -5734 297854 -4742
rect 300954 302614 301574 336000
rect 300954 302058 300986 302614
rect 301542 302058 301574 302614
rect 300954 266614 301574 302058
rect 300954 266058 300986 266614
rect 301542 266058 301574 266614
rect 300954 230614 301574 266058
rect 300954 230058 300986 230614
rect 301542 230058 301574 230614
rect 300954 194614 301574 230058
rect 300954 194058 300986 194614
rect 301542 194058 301574 194614
rect 300954 158614 301574 194058
rect 300954 158058 300986 158614
rect 301542 158058 301574 158614
rect 300954 122614 301574 158058
rect 300954 122058 300986 122614
rect 301542 122058 301574 122614
rect 300954 86614 301574 122058
rect 300954 86058 300986 86614
rect 301542 86058 301574 86614
rect 300954 50614 301574 86058
rect 300954 50058 300986 50614
rect 301542 50058 301574 50614
rect 300954 14614 301574 50058
rect 300954 14058 300986 14614
rect 301542 14058 301574 14614
rect 282954 -7622 282986 -7066
rect 283542 -7622 283574 -7066
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 309454 308414 336000
rect 307794 308898 307826 309454
rect 308382 308898 308414 309454
rect 307794 273454 308414 308898
rect 307794 272898 307826 273454
rect 308382 272898 308414 273454
rect 307794 237454 308414 272898
rect 307794 236898 307826 237454
rect 308382 236898 308414 237454
rect 307794 201454 308414 236898
rect 307794 200898 307826 201454
rect 308382 200898 308414 201454
rect 307794 165454 308414 200898
rect 307794 164898 307826 165454
rect 308382 164898 308414 165454
rect 307794 129454 308414 164898
rect 307794 128898 307826 129454
rect 308382 128898 308414 129454
rect 307794 93454 308414 128898
rect 307794 92898 307826 93454
rect 308382 92898 308414 93454
rect 307794 57454 308414 92898
rect 307794 56898 307826 57454
rect 308382 56898 308414 57454
rect 307794 21454 308414 56898
rect 307794 20898 307826 21454
rect 308382 20898 308414 21454
rect 307794 -1306 308414 20898
rect 307794 -1862 307826 -1306
rect 308382 -1862 308414 -1306
rect 307794 -1894 308414 -1862
rect 311514 313174 312134 336000
rect 311514 312618 311546 313174
rect 312102 312618 312134 313174
rect 311514 277174 312134 312618
rect 311514 276618 311546 277174
rect 312102 276618 312134 277174
rect 311514 241174 312134 276618
rect 311514 240618 311546 241174
rect 312102 240618 312134 241174
rect 311514 205174 312134 240618
rect 311514 204618 311546 205174
rect 312102 204618 312134 205174
rect 311514 169174 312134 204618
rect 311514 168618 311546 169174
rect 312102 168618 312134 169174
rect 311514 133174 312134 168618
rect 311514 132618 311546 133174
rect 312102 132618 312134 133174
rect 311514 97174 312134 132618
rect 311514 96618 311546 97174
rect 312102 96618 312134 97174
rect 311514 61174 312134 96618
rect 311514 60618 311546 61174
rect 312102 60618 312134 61174
rect 311514 25174 312134 60618
rect 311514 24618 311546 25174
rect 312102 24618 312134 25174
rect 311514 -3226 312134 24618
rect 311514 -3782 311546 -3226
rect 312102 -3782 312134 -3226
rect 311514 -3814 312134 -3782
rect 315234 316894 315854 336000
rect 315234 316338 315266 316894
rect 315822 316338 315854 316894
rect 315234 280894 315854 316338
rect 315234 280338 315266 280894
rect 315822 280338 315854 280894
rect 315234 244894 315854 280338
rect 315234 244338 315266 244894
rect 315822 244338 315854 244894
rect 315234 208894 315854 244338
rect 315234 208338 315266 208894
rect 315822 208338 315854 208894
rect 315234 172894 315854 208338
rect 315234 172338 315266 172894
rect 315822 172338 315854 172894
rect 315234 136894 315854 172338
rect 315234 136338 315266 136894
rect 315822 136338 315854 136894
rect 315234 100894 315854 136338
rect 315234 100338 315266 100894
rect 315822 100338 315854 100894
rect 315234 64894 315854 100338
rect 315234 64338 315266 64894
rect 315822 64338 315854 64894
rect 315234 28894 315854 64338
rect 315234 28338 315266 28894
rect 315822 28338 315854 28894
rect 315234 -5146 315854 28338
rect 315234 -5702 315266 -5146
rect 315822 -5702 315854 -5146
rect 315234 -5734 315854 -5702
rect 318954 320614 319574 336000
rect 318954 320058 318986 320614
rect 319542 320058 319574 320614
rect 318954 284614 319574 320058
rect 318954 284058 318986 284614
rect 319542 284058 319574 284614
rect 318954 248614 319574 284058
rect 318954 248058 318986 248614
rect 319542 248058 319574 248614
rect 318954 212614 319574 248058
rect 318954 212058 318986 212614
rect 319542 212058 319574 212614
rect 318954 176614 319574 212058
rect 318954 176058 318986 176614
rect 319542 176058 319574 176614
rect 318954 140614 319574 176058
rect 318954 140058 318986 140614
rect 319542 140058 319574 140614
rect 318954 104614 319574 140058
rect 318954 104058 318986 104614
rect 319542 104058 319574 104614
rect 318954 68614 319574 104058
rect 318954 68058 318986 68614
rect 319542 68058 319574 68614
rect 318954 32614 319574 68058
rect 318954 32058 318986 32614
rect 319542 32058 319574 32614
rect 300954 -6662 300986 -6106
rect 301542 -6662 301574 -6106
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 327454 326414 336000
rect 325794 326898 325826 327454
rect 326382 326898 326414 327454
rect 325794 291454 326414 326898
rect 325794 290898 325826 291454
rect 326382 290898 326414 291454
rect 325794 255454 326414 290898
rect 325794 254898 325826 255454
rect 326382 254898 326414 255454
rect 325794 219454 326414 254898
rect 325794 218898 325826 219454
rect 326382 218898 326414 219454
rect 325794 183454 326414 218898
rect 325794 182898 325826 183454
rect 326382 182898 326414 183454
rect 325794 147454 326414 182898
rect 325794 146898 325826 147454
rect 326382 146898 326414 147454
rect 325794 111454 326414 146898
rect 325794 110898 325826 111454
rect 326382 110898 326414 111454
rect 325794 75454 326414 110898
rect 325794 74898 325826 75454
rect 326382 74898 326414 75454
rect 325794 39454 326414 74898
rect 325794 38898 325826 39454
rect 326382 38898 326414 39454
rect 325794 3454 326414 38898
rect 325794 2898 325826 3454
rect 326382 2898 326414 3454
rect 325794 -346 326414 2898
rect 325794 -902 325826 -346
rect 326382 -902 326414 -346
rect 325794 -1894 326414 -902
rect 329514 331174 330134 336000
rect 329514 330618 329546 331174
rect 330102 330618 330134 331174
rect 329514 295174 330134 330618
rect 329514 294618 329546 295174
rect 330102 294618 330134 295174
rect 329514 259174 330134 294618
rect 329514 258618 329546 259174
rect 330102 258618 330134 259174
rect 329514 223174 330134 258618
rect 329514 222618 329546 223174
rect 330102 222618 330134 223174
rect 329514 187174 330134 222618
rect 329514 186618 329546 187174
rect 330102 186618 330134 187174
rect 329514 151174 330134 186618
rect 329514 150618 329546 151174
rect 330102 150618 330134 151174
rect 329514 115174 330134 150618
rect 329514 114618 329546 115174
rect 330102 114618 330134 115174
rect 329514 79174 330134 114618
rect 329514 78618 329546 79174
rect 330102 78618 330134 79174
rect 329514 43174 330134 78618
rect 329514 42618 329546 43174
rect 330102 42618 330134 43174
rect 329514 7174 330134 42618
rect 329514 6618 329546 7174
rect 330102 6618 330134 7174
rect 329514 -2266 330134 6618
rect 329514 -2822 329546 -2266
rect 330102 -2822 330134 -2266
rect 329514 -3814 330134 -2822
rect 333234 334894 333854 336000
rect 333234 334338 333266 334894
rect 333822 334338 333854 334894
rect 333234 298894 333854 334338
rect 333234 298338 333266 298894
rect 333822 298338 333854 298894
rect 333234 262894 333854 298338
rect 333234 262338 333266 262894
rect 333822 262338 333854 262894
rect 333234 226894 333854 262338
rect 333234 226338 333266 226894
rect 333822 226338 333854 226894
rect 333234 190894 333854 226338
rect 333234 190338 333266 190894
rect 333822 190338 333854 190894
rect 333234 154894 333854 190338
rect 333234 154338 333266 154894
rect 333822 154338 333854 154894
rect 333234 118894 333854 154338
rect 333234 118338 333266 118894
rect 333822 118338 333854 118894
rect 333234 82894 333854 118338
rect 333234 82338 333266 82894
rect 333822 82338 333854 82894
rect 333234 46894 333854 82338
rect 333234 46338 333266 46894
rect 333822 46338 333854 46894
rect 333234 10894 333854 46338
rect 333234 10338 333266 10894
rect 333822 10338 333854 10894
rect 333234 -4186 333854 10338
rect 333234 -4742 333266 -4186
rect 333822 -4742 333854 -4186
rect 333234 -5734 333854 -4742
rect 336954 302614 337574 336000
rect 336954 302058 336986 302614
rect 337542 302058 337574 302614
rect 336954 266614 337574 302058
rect 336954 266058 336986 266614
rect 337542 266058 337574 266614
rect 336954 230614 337574 266058
rect 336954 230058 336986 230614
rect 337542 230058 337574 230614
rect 336954 194614 337574 230058
rect 336954 194058 336986 194614
rect 337542 194058 337574 194614
rect 336954 158614 337574 194058
rect 336954 158058 336986 158614
rect 337542 158058 337574 158614
rect 336954 122614 337574 158058
rect 336954 122058 336986 122614
rect 337542 122058 337574 122614
rect 336954 86614 337574 122058
rect 336954 86058 336986 86614
rect 337542 86058 337574 86614
rect 336954 50614 337574 86058
rect 336954 50058 336986 50614
rect 337542 50058 337574 50614
rect 336954 14614 337574 50058
rect 336954 14058 336986 14614
rect 337542 14058 337574 14614
rect 318954 -7622 318986 -7066
rect 319542 -7622 319574 -7066
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 309454 344414 336000
rect 343794 308898 343826 309454
rect 344382 308898 344414 309454
rect 343794 273454 344414 308898
rect 343794 272898 343826 273454
rect 344382 272898 344414 273454
rect 343794 237454 344414 272898
rect 343794 236898 343826 237454
rect 344382 236898 344414 237454
rect 343794 201454 344414 236898
rect 343794 200898 343826 201454
rect 344382 200898 344414 201454
rect 343794 165454 344414 200898
rect 343794 164898 343826 165454
rect 344382 164898 344414 165454
rect 343794 129454 344414 164898
rect 343794 128898 343826 129454
rect 344382 128898 344414 129454
rect 343794 93454 344414 128898
rect 343794 92898 343826 93454
rect 344382 92898 344414 93454
rect 343794 57454 344414 92898
rect 343794 56898 343826 57454
rect 344382 56898 344414 57454
rect 343794 21454 344414 56898
rect 343794 20898 343826 21454
rect 344382 20898 344414 21454
rect 343794 -1306 344414 20898
rect 343794 -1862 343826 -1306
rect 344382 -1862 344414 -1306
rect 343794 -1894 344414 -1862
rect 347514 313174 348134 336000
rect 347514 312618 347546 313174
rect 348102 312618 348134 313174
rect 347514 277174 348134 312618
rect 347514 276618 347546 277174
rect 348102 276618 348134 277174
rect 347514 241174 348134 276618
rect 347514 240618 347546 241174
rect 348102 240618 348134 241174
rect 347514 205174 348134 240618
rect 347514 204618 347546 205174
rect 348102 204618 348134 205174
rect 347514 169174 348134 204618
rect 347514 168618 347546 169174
rect 348102 168618 348134 169174
rect 347514 133174 348134 168618
rect 347514 132618 347546 133174
rect 348102 132618 348134 133174
rect 347514 97174 348134 132618
rect 347514 96618 347546 97174
rect 348102 96618 348134 97174
rect 347514 61174 348134 96618
rect 347514 60618 347546 61174
rect 348102 60618 348134 61174
rect 347514 25174 348134 60618
rect 347514 24618 347546 25174
rect 348102 24618 348134 25174
rect 347514 -3226 348134 24618
rect 347514 -3782 347546 -3226
rect 348102 -3782 348134 -3226
rect 347514 -3814 348134 -3782
rect 351234 316894 351854 336000
rect 351234 316338 351266 316894
rect 351822 316338 351854 316894
rect 351234 280894 351854 316338
rect 351234 280338 351266 280894
rect 351822 280338 351854 280894
rect 351234 244894 351854 280338
rect 351234 244338 351266 244894
rect 351822 244338 351854 244894
rect 351234 208894 351854 244338
rect 351234 208338 351266 208894
rect 351822 208338 351854 208894
rect 351234 172894 351854 208338
rect 351234 172338 351266 172894
rect 351822 172338 351854 172894
rect 351234 136894 351854 172338
rect 351234 136338 351266 136894
rect 351822 136338 351854 136894
rect 351234 100894 351854 136338
rect 351234 100338 351266 100894
rect 351822 100338 351854 100894
rect 351234 64894 351854 100338
rect 351234 64338 351266 64894
rect 351822 64338 351854 64894
rect 351234 28894 351854 64338
rect 351234 28338 351266 28894
rect 351822 28338 351854 28894
rect 351234 -5146 351854 28338
rect 351234 -5702 351266 -5146
rect 351822 -5702 351854 -5146
rect 351234 -5734 351854 -5702
rect 354954 320614 355574 336000
rect 354954 320058 354986 320614
rect 355542 320058 355574 320614
rect 354954 284614 355574 320058
rect 354954 284058 354986 284614
rect 355542 284058 355574 284614
rect 354954 248614 355574 284058
rect 354954 248058 354986 248614
rect 355542 248058 355574 248614
rect 354954 212614 355574 248058
rect 354954 212058 354986 212614
rect 355542 212058 355574 212614
rect 354954 176614 355574 212058
rect 354954 176058 354986 176614
rect 355542 176058 355574 176614
rect 354954 140614 355574 176058
rect 354954 140058 354986 140614
rect 355542 140058 355574 140614
rect 354954 104614 355574 140058
rect 354954 104058 354986 104614
rect 355542 104058 355574 104614
rect 354954 68614 355574 104058
rect 354954 68058 354986 68614
rect 355542 68058 355574 68614
rect 354954 32614 355574 68058
rect 354954 32058 354986 32614
rect 355542 32058 355574 32614
rect 336954 -6662 336986 -6106
rect 337542 -6662 337574 -6106
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 327454 362414 336000
rect 361794 326898 361826 327454
rect 362382 326898 362414 327454
rect 361794 291454 362414 326898
rect 361794 290898 361826 291454
rect 362382 290898 362414 291454
rect 361794 255454 362414 290898
rect 361794 254898 361826 255454
rect 362382 254898 362414 255454
rect 361794 219454 362414 254898
rect 361794 218898 361826 219454
rect 362382 218898 362414 219454
rect 361794 183454 362414 218898
rect 361794 182898 361826 183454
rect 362382 182898 362414 183454
rect 361794 147454 362414 182898
rect 361794 146898 361826 147454
rect 362382 146898 362414 147454
rect 361794 111454 362414 146898
rect 361794 110898 361826 111454
rect 362382 110898 362414 111454
rect 361794 75454 362414 110898
rect 361794 74898 361826 75454
rect 362382 74898 362414 75454
rect 361794 39454 362414 74898
rect 361794 38898 361826 39454
rect 362382 38898 362414 39454
rect 361794 3454 362414 38898
rect 361794 2898 361826 3454
rect 362382 2898 362414 3454
rect 361794 -346 362414 2898
rect 361794 -902 361826 -346
rect 362382 -902 362414 -346
rect 361794 -1894 362414 -902
rect 365514 331174 366134 336000
rect 365514 330618 365546 331174
rect 366102 330618 366134 331174
rect 365514 295174 366134 330618
rect 365514 294618 365546 295174
rect 366102 294618 366134 295174
rect 365514 259174 366134 294618
rect 365514 258618 365546 259174
rect 366102 258618 366134 259174
rect 365514 223174 366134 258618
rect 365514 222618 365546 223174
rect 366102 222618 366134 223174
rect 365514 187174 366134 222618
rect 365514 186618 365546 187174
rect 366102 186618 366134 187174
rect 365514 151174 366134 186618
rect 365514 150618 365546 151174
rect 366102 150618 366134 151174
rect 365514 115174 366134 150618
rect 365514 114618 365546 115174
rect 366102 114618 366134 115174
rect 365514 79174 366134 114618
rect 365514 78618 365546 79174
rect 366102 78618 366134 79174
rect 365514 43174 366134 78618
rect 365514 42618 365546 43174
rect 366102 42618 366134 43174
rect 365514 7174 366134 42618
rect 365514 6618 365546 7174
rect 366102 6618 366134 7174
rect 365514 -2266 366134 6618
rect 365514 -2822 365546 -2266
rect 366102 -2822 366134 -2266
rect 365514 -3814 366134 -2822
rect 369234 334894 369854 336000
rect 369234 334338 369266 334894
rect 369822 334338 369854 334894
rect 369234 298894 369854 334338
rect 369234 298338 369266 298894
rect 369822 298338 369854 298894
rect 369234 262894 369854 298338
rect 369234 262338 369266 262894
rect 369822 262338 369854 262894
rect 369234 226894 369854 262338
rect 369234 226338 369266 226894
rect 369822 226338 369854 226894
rect 369234 190894 369854 226338
rect 369234 190338 369266 190894
rect 369822 190338 369854 190894
rect 369234 154894 369854 190338
rect 369234 154338 369266 154894
rect 369822 154338 369854 154894
rect 369234 118894 369854 154338
rect 369234 118338 369266 118894
rect 369822 118338 369854 118894
rect 369234 82894 369854 118338
rect 369234 82338 369266 82894
rect 369822 82338 369854 82894
rect 369234 46894 369854 82338
rect 369234 46338 369266 46894
rect 369822 46338 369854 46894
rect 369234 10894 369854 46338
rect 369234 10338 369266 10894
rect 369822 10338 369854 10894
rect 369234 -4186 369854 10338
rect 369234 -4742 369266 -4186
rect 369822 -4742 369854 -4186
rect 369234 -5734 369854 -4742
rect 372954 302614 373574 336000
rect 372954 302058 372986 302614
rect 373542 302058 373574 302614
rect 372954 266614 373574 302058
rect 372954 266058 372986 266614
rect 373542 266058 373574 266614
rect 372954 230614 373574 266058
rect 372954 230058 372986 230614
rect 373542 230058 373574 230614
rect 372954 194614 373574 230058
rect 372954 194058 372986 194614
rect 373542 194058 373574 194614
rect 372954 158614 373574 194058
rect 372954 158058 372986 158614
rect 373542 158058 373574 158614
rect 372954 122614 373574 158058
rect 372954 122058 372986 122614
rect 373542 122058 373574 122614
rect 372954 86614 373574 122058
rect 372954 86058 372986 86614
rect 373542 86058 373574 86614
rect 372954 50614 373574 86058
rect 372954 50058 372986 50614
rect 373542 50058 373574 50614
rect 372954 14614 373574 50058
rect 372954 14058 372986 14614
rect 373542 14058 373574 14614
rect 354954 -7622 354986 -7066
rect 355542 -7622 355574 -7066
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 309454 380414 336000
rect 379794 308898 379826 309454
rect 380382 308898 380414 309454
rect 379794 273454 380414 308898
rect 379794 272898 379826 273454
rect 380382 272898 380414 273454
rect 379794 237454 380414 272898
rect 379794 236898 379826 237454
rect 380382 236898 380414 237454
rect 379794 201454 380414 236898
rect 379794 200898 379826 201454
rect 380382 200898 380414 201454
rect 379794 165454 380414 200898
rect 379794 164898 379826 165454
rect 380382 164898 380414 165454
rect 379794 129454 380414 164898
rect 379794 128898 379826 129454
rect 380382 128898 380414 129454
rect 379794 93454 380414 128898
rect 379794 92898 379826 93454
rect 380382 92898 380414 93454
rect 379794 57454 380414 92898
rect 379794 56898 379826 57454
rect 380382 56898 380414 57454
rect 379794 21454 380414 56898
rect 379794 20898 379826 21454
rect 380382 20898 380414 21454
rect 379794 -1306 380414 20898
rect 379794 -1862 379826 -1306
rect 380382 -1862 380414 -1306
rect 379794 -1894 380414 -1862
rect 383514 313174 384134 336000
rect 383514 312618 383546 313174
rect 384102 312618 384134 313174
rect 383514 277174 384134 312618
rect 383514 276618 383546 277174
rect 384102 276618 384134 277174
rect 383514 241174 384134 276618
rect 383514 240618 383546 241174
rect 384102 240618 384134 241174
rect 383514 205174 384134 240618
rect 383514 204618 383546 205174
rect 384102 204618 384134 205174
rect 383514 169174 384134 204618
rect 383514 168618 383546 169174
rect 384102 168618 384134 169174
rect 383514 133174 384134 168618
rect 383514 132618 383546 133174
rect 384102 132618 384134 133174
rect 383514 97174 384134 132618
rect 383514 96618 383546 97174
rect 384102 96618 384134 97174
rect 383514 61174 384134 96618
rect 383514 60618 383546 61174
rect 384102 60618 384134 61174
rect 383514 25174 384134 60618
rect 383514 24618 383546 25174
rect 384102 24618 384134 25174
rect 383514 -3226 384134 24618
rect 383514 -3782 383546 -3226
rect 384102 -3782 384134 -3226
rect 383514 -3814 384134 -3782
rect 387234 316894 387854 336000
rect 387234 316338 387266 316894
rect 387822 316338 387854 316894
rect 387234 280894 387854 316338
rect 387234 280338 387266 280894
rect 387822 280338 387854 280894
rect 387234 244894 387854 280338
rect 387234 244338 387266 244894
rect 387822 244338 387854 244894
rect 387234 208894 387854 244338
rect 387234 208338 387266 208894
rect 387822 208338 387854 208894
rect 387234 172894 387854 208338
rect 387234 172338 387266 172894
rect 387822 172338 387854 172894
rect 387234 136894 387854 172338
rect 387234 136338 387266 136894
rect 387822 136338 387854 136894
rect 387234 100894 387854 136338
rect 387234 100338 387266 100894
rect 387822 100338 387854 100894
rect 387234 64894 387854 100338
rect 387234 64338 387266 64894
rect 387822 64338 387854 64894
rect 387234 28894 387854 64338
rect 387234 28338 387266 28894
rect 387822 28338 387854 28894
rect 387234 -5146 387854 28338
rect 387234 -5702 387266 -5146
rect 387822 -5702 387854 -5146
rect 387234 -5734 387854 -5702
rect 390954 320614 391574 336000
rect 390954 320058 390986 320614
rect 391542 320058 391574 320614
rect 390954 284614 391574 320058
rect 390954 284058 390986 284614
rect 391542 284058 391574 284614
rect 390954 248614 391574 284058
rect 390954 248058 390986 248614
rect 391542 248058 391574 248614
rect 390954 212614 391574 248058
rect 390954 212058 390986 212614
rect 391542 212058 391574 212614
rect 390954 176614 391574 212058
rect 390954 176058 390986 176614
rect 391542 176058 391574 176614
rect 390954 140614 391574 176058
rect 390954 140058 390986 140614
rect 391542 140058 391574 140614
rect 390954 104614 391574 140058
rect 390954 104058 390986 104614
rect 391542 104058 391574 104614
rect 390954 68614 391574 104058
rect 390954 68058 390986 68614
rect 391542 68058 391574 68614
rect 390954 32614 391574 68058
rect 390954 32058 390986 32614
rect 391542 32058 391574 32614
rect 372954 -6662 372986 -6106
rect 373542 -6662 373574 -6106
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 327454 398414 336000
rect 397794 326898 397826 327454
rect 398382 326898 398414 327454
rect 397794 291454 398414 326898
rect 397794 290898 397826 291454
rect 398382 290898 398414 291454
rect 397794 255454 398414 290898
rect 397794 254898 397826 255454
rect 398382 254898 398414 255454
rect 397794 219454 398414 254898
rect 397794 218898 397826 219454
rect 398382 218898 398414 219454
rect 397794 183454 398414 218898
rect 397794 182898 397826 183454
rect 398382 182898 398414 183454
rect 397794 147454 398414 182898
rect 397794 146898 397826 147454
rect 398382 146898 398414 147454
rect 397794 111454 398414 146898
rect 397794 110898 397826 111454
rect 398382 110898 398414 111454
rect 397794 75454 398414 110898
rect 397794 74898 397826 75454
rect 398382 74898 398414 75454
rect 397794 39454 398414 74898
rect 397794 38898 397826 39454
rect 398382 38898 398414 39454
rect 397794 3454 398414 38898
rect 397794 2898 397826 3454
rect 398382 2898 398414 3454
rect 397794 -346 398414 2898
rect 397794 -902 397826 -346
rect 398382 -902 398414 -346
rect 397794 -1894 398414 -902
rect 401514 331174 402134 336000
rect 401514 330618 401546 331174
rect 402102 330618 402134 331174
rect 401514 295174 402134 330618
rect 401514 294618 401546 295174
rect 402102 294618 402134 295174
rect 401514 259174 402134 294618
rect 401514 258618 401546 259174
rect 402102 258618 402134 259174
rect 401514 223174 402134 258618
rect 401514 222618 401546 223174
rect 402102 222618 402134 223174
rect 401514 187174 402134 222618
rect 401514 186618 401546 187174
rect 402102 186618 402134 187174
rect 401514 151174 402134 186618
rect 401514 150618 401546 151174
rect 402102 150618 402134 151174
rect 401514 115174 402134 150618
rect 401514 114618 401546 115174
rect 402102 114618 402134 115174
rect 401514 79174 402134 114618
rect 401514 78618 401546 79174
rect 402102 78618 402134 79174
rect 401514 43174 402134 78618
rect 401514 42618 401546 43174
rect 402102 42618 402134 43174
rect 401514 7174 402134 42618
rect 401514 6618 401546 7174
rect 402102 6618 402134 7174
rect 401514 -2266 402134 6618
rect 401514 -2822 401546 -2266
rect 402102 -2822 402134 -2266
rect 401514 -3814 402134 -2822
rect 405234 334894 405854 336000
rect 405234 334338 405266 334894
rect 405822 334338 405854 334894
rect 405234 298894 405854 334338
rect 405234 298338 405266 298894
rect 405822 298338 405854 298894
rect 405234 262894 405854 298338
rect 405234 262338 405266 262894
rect 405822 262338 405854 262894
rect 405234 226894 405854 262338
rect 405234 226338 405266 226894
rect 405822 226338 405854 226894
rect 405234 190894 405854 226338
rect 405234 190338 405266 190894
rect 405822 190338 405854 190894
rect 405234 154894 405854 190338
rect 405234 154338 405266 154894
rect 405822 154338 405854 154894
rect 405234 118894 405854 154338
rect 405234 118338 405266 118894
rect 405822 118338 405854 118894
rect 405234 82894 405854 118338
rect 405234 82338 405266 82894
rect 405822 82338 405854 82894
rect 405234 46894 405854 82338
rect 405234 46338 405266 46894
rect 405822 46338 405854 46894
rect 405234 10894 405854 46338
rect 405234 10338 405266 10894
rect 405822 10338 405854 10894
rect 405234 -4186 405854 10338
rect 405234 -4742 405266 -4186
rect 405822 -4742 405854 -4186
rect 405234 -5734 405854 -4742
rect 408954 302614 409574 336000
rect 408954 302058 408986 302614
rect 409542 302058 409574 302614
rect 408954 266614 409574 302058
rect 408954 266058 408986 266614
rect 409542 266058 409574 266614
rect 408954 230614 409574 266058
rect 408954 230058 408986 230614
rect 409542 230058 409574 230614
rect 408954 194614 409574 230058
rect 408954 194058 408986 194614
rect 409542 194058 409574 194614
rect 408954 158614 409574 194058
rect 408954 158058 408986 158614
rect 409542 158058 409574 158614
rect 408954 122614 409574 158058
rect 408954 122058 408986 122614
rect 409542 122058 409574 122614
rect 408954 86614 409574 122058
rect 408954 86058 408986 86614
rect 409542 86058 409574 86614
rect 408954 50614 409574 86058
rect 408954 50058 408986 50614
rect 409542 50058 409574 50614
rect 408954 14614 409574 50058
rect 408954 14058 408986 14614
rect 409542 14058 409574 14614
rect 390954 -7622 390986 -7066
rect 391542 -7622 391574 -7066
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 309454 416414 336000
rect 415794 308898 415826 309454
rect 416382 308898 416414 309454
rect 415794 273454 416414 308898
rect 415794 272898 415826 273454
rect 416382 272898 416414 273454
rect 415794 237454 416414 272898
rect 415794 236898 415826 237454
rect 416382 236898 416414 237454
rect 415794 201454 416414 236898
rect 415794 200898 415826 201454
rect 416382 200898 416414 201454
rect 415794 165454 416414 200898
rect 415794 164898 415826 165454
rect 416382 164898 416414 165454
rect 415794 129454 416414 164898
rect 415794 128898 415826 129454
rect 416382 128898 416414 129454
rect 415794 93454 416414 128898
rect 415794 92898 415826 93454
rect 416382 92898 416414 93454
rect 415794 57454 416414 92898
rect 415794 56898 415826 57454
rect 416382 56898 416414 57454
rect 415794 21454 416414 56898
rect 415794 20898 415826 21454
rect 416382 20898 416414 21454
rect 415794 -1306 416414 20898
rect 415794 -1862 415826 -1306
rect 416382 -1862 416414 -1306
rect 415794 -1894 416414 -1862
rect 419514 313174 420134 336000
rect 419514 312618 419546 313174
rect 420102 312618 420134 313174
rect 419514 277174 420134 312618
rect 419514 276618 419546 277174
rect 420102 276618 420134 277174
rect 419514 241174 420134 276618
rect 419514 240618 419546 241174
rect 420102 240618 420134 241174
rect 419514 205174 420134 240618
rect 419514 204618 419546 205174
rect 420102 204618 420134 205174
rect 419514 169174 420134 204618
rect 419514 168618 419546 169174
rect 420102 168618 420134 169174
rect 419514 133174 420134 168618
rect 419514 132618 419546 133174
rect 420102 132618 420134 133174
rect 419514 97174 420134 132618
rect 419514 96618 419546 97174
rect 420102 96618 420134 97174
rect 419514 61174 420134 96618
rect 419514 60618 419546 61174
rect 420102 60618 420134 61174
rect 419514 25174 420134 60618
rect 419514 24618 419546 25174
rect 420102 24618 420134 25174
rect 419514 -3226 420134 24618
rect 419514 -3782 419546 -3226
rect 420102 -3782 420134 -3226
rect 419514 -3814 420134 -3782
rect 423234 316894 423854 336000
rect 423234 316338 423266 316894
rect 423822 316338 423854 316894
rect 423234 280894 423854 316338
rect 423234 280338 423266 280894
rect 423822 280338 423854 280894
rect 423234 244894 423854 280338
rect 423234 244338 423266 244894
rect 423822 244338 423854 244894
rect 423234 208894 423854 244338
rect 423234 208338 423266 208894
rect 423822 208338 423854 208894
rect 423234 172894 423854 208338
rect 423234 172338 423266 172894
rect 423822 172338 423854 172894
rect 423234 136894 423854 172338
rect 423234 136338 423266 136894
rect 423822 136338 423854 136894
rect 423234 100894 423854 136338
rect 423234 100338 423266 100894
rect 423822 100338 423854 100894
rect 423234 64894 423854 100338
rect 423998 96661 424058 497387
rect 423995 96660 424061 96661
rect 423995 96596 423996 96660
rect 424060 96596 424061 96660
rect 423995 96595 424061 96596
rect 425102 70413 425162 497387
rect 425099 70412 425165 70413
rect 425099 70348 425100 70412
rect 425164 70348 425165 70412
rect 425099 70347 425165 70348
rect 423234 64338 423266 64894
rect 423822 64338 423854 64894
rect 423234 28894 423854 64338
rect 426390 44301 426450 497387
rect 426954 320614 427574 336000
rect 426954 320058 426986 320614
rect 427542 320058 427574 320614
rect 426954 284614 427574 320058
rect 426954 284058 426986 284614
rect 427542 284058 427574 284614
rect 426954 248614 427574 284058
rect 426954 248058 426986 248614
rect 427542 248058 427574 248614
rect 426954 212614 427574 248058
rect 426954 212058 426986 212614
rect 427542 212058 427574 212614
rect 426954 176614 427574 212058
rect 426954 176058 426986 176614
rect 427542 176058 427574 176614
rect 426954 140614 427574 176058
rect 426954 140058 426986 140614
rect 427542 140058 427574 140614
rect 426954 104614 427574 140058
rect 426954 104058 426986 104614
rect 427542 104058 427574 104614
rect 426954 68614 427574 104058
rect 426954 68058 426986 68614
rect 427542 68058 427574 68614
rect 426387 44300 426453 44301
rect 426387 44236 426388 44300
rect 426452 44236 426453 44300
rect 426387 44235 426453 44236
rect 423234 28338 423266 28894
rect 423822 28338 423854 28894
rect 423234 -5146 423854 28338
rect 423234 -5702 423266 -5146
rect 423822 -5702 423854 -5146
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 68058
rect 427862 58037 427922 497387
rect 427859 58036 427925 58037
rect 427859 57972 427860 58036
rect 427924 57972 427925 58036
rect 427859 57971 427925 57972
rect 426954 32058 426986 32614
rect 427542 32058 427574 32614
rect 408954 -6662 408986 -6106
rect 409542 -6662 409574 -6106
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 429150 31789 429210 497387
rect 429147 31788 429213 31789
rect 429147 31724 429148 31788
rect 429212 31724 429213 31788
rect 429147 31723 429213 31724
rect 433382 19413 433442 497387
rect 437514 475174 438134 510618
rect 437514 474618 437546 475174
rect 438102 474618 438134 475174
rect 437514 439174 438134 474618
rect 437514 438618 437546 439174
rect 438102 438618 438134 439174
rect 437514 403174 438134 438618
rect 437514 402618 437546 403174
rect 438102 402618 438134 403174
rect 437514 367174 438134 402618
rect 437514 366618 437546 367174
rect 438102 366618 438134 367174
rect 433794 327454 434414 336000
rect 433794 326898 433826 327454
rect 434382 326898 434414 327454
rect 433794 291454 434414 326898
rect 433794 290898 433826 291454
rect 434382 290898 434414 291454
rect 433794 255454 434414 290898
rect 433794 254898 433826 255454
rect 434382 254898 434414 255454
rect 433794 219454 434414 254898
rect 433794 218898 433826 219454
rect 434382 218898 434414 219454
rect 433794 183454 434414 218898
rect 433794 182898 433826 183454
rect 434382 182898 434414 183454
rect 433794 147454 434414 182898
rect 433794 146898 433826 147454
rect 434382 146898 434414 147454
rect 433794 111454 434414 146898
rect 433794 110898 433826 111454
rect 434382 110898 434414 111454
rect 433794 75454 434414 110898
rect 433794 74898 433826 75454
rect 434382 74898 434414 75454
rect 433794 39454 434414 74898
rect 433794 38898 433826 39454
rect 434382 38898 434414 39454
rect 433379 19412 433445 19413
rect 433379 19348 433380 19412
rect 433444 19348 433445 19412
rect 433379 19347 433445 19348
rect 433794 3454 434414 38898
rect 433794 2898 433826 3454
rect 434382 2898 434414 3454
rect 433794 -346 434414 2898
rect 433794 -902 433826 -346
rect 434382 -902 434414 -346
rect 433794 -1894 434414 -902
rect 437514 331174 438134 366618
rect 437514 330618 437546 331174
rect 438102 330618 438134 331174
rect 437514 295174 438134 330618
rect 437514 294618 437546 295174
rect 438102 294618 438134 295174
rect 437514 259174 438134 294618
rect 437514 258618 437546 259174
rect 438102 258618 438134 259174
rect 437514 223174 438134 258618
rect 437514 222618 437546 223174
rect 438102 222618 438134 223174
rect 437514 187174 438134 222618
rect 437514 186618 437546 187174
rect 438102 186618 438134 187174
rect 437514 151174 438134 186618
rect 437514 150618 437546 151174
rect 438102 150618 438134 151174
rect 437514 115174 438134 150618
rect 437514 114618 437546 115174
rect 438102 114618 438134 115174
rect 437514 79174 438134 114618
rect 437514 78618 437546 79174
rect 438102 78618 438134 79174
rect 437514 43174 438134 78618
rect 437514 42618 437546 43174
rect 438102 42618 438134 43174
rect 437514 7174 438134 42618
rect 437514 6618 437546 7174
rect 438102 6618 438134 7174
rect 437514 -2266 438134 6618
rect 437514 -2822 437546 -2266
rect 438102 -2822 438134 -2266
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694338 441266 694894
rect 441822 694338 441854 694894
rect 441234 658894 441854 694338
rect 441234 658338 441266 658894
rect 441822 658338 441854 658894
rect 441234 622894 441854 658338
rect 441234 622338 441266 622894
rect 441822 622338 441854 622894
rect 441234 586894 441854 622338
rect 441234 586338 441266 586894
rect 441822 586338 441854 586894
rect 441234 550894 441854 586338
rect 441234 550338 441266 550894
rect 441822 550338 441854 550894
rect 441234 514894 441854 550338
rect 441234 514338 441266 514894
rect 441822 514338 441854 514894
rect 441234 478894 441854 514338
rect 441234 478338 441266 478894
rect 441822 478338 441854 478894
rect 441234 442894 441854 478338
rect 441234 442338 441266 442894
rect 441822 442338 441854 442894
rect 441234 406894 441854 442338
rect 441234 406338 441266 406894
rect 441822 406338 441854 406894
rect 441234 370894 441854 406338
rect 441234 370338 441266 370894
rect 441822 370338 441854 370894
rect 441234 334894 441854 370338
rect 441234 334338 441266 334894
rect 441822 334338 441854 334894
rect 441234 298894 441854 334338
rect 441234 298338 441266 298894
rect 441822 298338 441854 298894
rect 441234 262894 441854 298338
rect 441234 262338 441266 262894
rect 441822 262338 441854 262894
rect 441234 226894 441854 262338
rect 441234 226338 441266 226894
rect 441822 226338 441854 226894
rect 441234 190894 441854 226338
rect 441234 190338 441266 190894
rect 441822 190338 441854 190894
rect 441234 154894 441854 190338
rect 441234 154338 441266 154894
rect 441822 154338 441854 154894
rect 441234 118894 441854 154338
rect 441234 118338 441266 118894
rect 441822 118338 441854 118894
rect 441234 82894 441854 118338
rect 441234 82338 441266 82894
rect 441822 82338 441854 82894
rect 441234 46894 441854 82338
rect 441234 46338 441266 46894
rect 441822 46338 441854 46894
rect 441234 10894 441854 46338
rect 441234 10338 441266 10894
rect 441822 10338 441854 10894
rect 441234 -4186 441854 10338
rect 441234 -4742 441266 -4186
rect 441822 -4742 441854 -4186
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711002 462986 711558
rect 463542 711002 463574 711558
rect 459234 709638 459854 709670
rect 459234 709082 459266 709638
rect 459822 709082 459854 709638
rect 455514 707718 456134 707750
rect 455514 707162 455546 707718
rect 456102 707162 456134 707718
rect 444954 698058 444986 698614
rect 445542 698058 445574 698614
rect 444954 662614 445574 698058
rect 444954 662058 444986 662614
rect 445542 662058 445574 662614
rect 444954 626614 445574 662058
rect 444954 626058 444986 626614
rect 445542 626058 445574 626614
rect 444954 590614 445574 626058
rect 444954 590058 444986 590614
rect 445542 590058 445574 590614
rect 444954 554614 445574 590058
rect 444954 554058 444986 554614
rect 445542 554058 445574 554614
rect 444954 518614 445574 554058
rect 444954 518058 444986 518614
rect 445542 518058 445574 518614
rect 444954 482614 445574 518058
rect 444954 482058 444986 482614
rect 445542 482058 445574 482614
rect 444954 446614 445574 482058
rect 444954 446058 444986 446614
rect 445542 446058 445574 446614
rect 444954 410614 445574 446058
rect 444954 410058 444986 410614
rect 445542 410058 445574 410614
rect 444954 374614 445574 410058
rect 444954 374058 444986 374614
rect 445542 374058 445574 374614
rect 444954 338614 445574 374058
rect 444954 338058 444986 338614
rect 445542 338058 445574 338614
rect 444954 302614 445574 338058
rect 444954 302058 444986 302614
rect 445542 302058 445574 302614
rect 444954 266614 445574 302058
rect 444954 266058 444986 266614
rect 445542 266058 445574 266614
rect 444954 230614 445574 266058
rect 444954 230058 444986 230614
rect 445542 230058 445574 230614
rect 444954 194614 445574 230058
rect 444954 194058 444986 194614
rect 445542 194058 445574 194614
rect 444954 158614 445574 194058
rect 444954 158058 444986 158614
rect 445542 158058 445574 158614
rect 444954 122614 445574 158058
rect 444954 122058 444986 122614
rect 445542 122058 445574 122614
rect 444954 86614 445574 122058
rect 444954 86058 444986 86614
rect 445542 86058 445574 86614
rect 444954 50614 445574 86058
rect 444954 50058 444986 50614
rect 445542 50058 445574 50614
rect 444954 14614 445574 50058
rect 444954 14058 444986 14614
rect 445542 14058 445574 14614
rect 426954 -7622 426986 -7066
rect 427542 -7622 427574 -7066
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705242 451826 705798
rect 452382 705242 452414 705798
rect 451794 669454 452414 705242
rect 451794 668898 451826 669454
rect 452382 668898 452414 669454
rect 451794 633454 452414 668898
rect 451794 632898 451826 633454
rect 452382 632898 452414 633454
rect 451794 597454 452414 632898
rect 451794 596898 451826 597454
rect 452382 596898 452414 597454
rect 451794 561454 452414 596898
rect 451794 560898 451826 561454
rect 452382 560898 452414 561454
rect 451794 525454 452414 560898
rect 451794 524898 451826 525454
rect 452382 524898 452414 525454
rect 451794 489454 452414 524898
rect 451794 488898 451826 489454
rect 452382 488898 452414 489454
rect 451794 453454 452414 488898
rect 451794 452898 451826 453454
rect 452382 452898 452414 453454
rect 451794 417454 452414 452898
rect 451794 416898 451826 417454
rect 452382 416898 452414 417454
rect 451794 381454 452414 416898
rect 451794 380898 451826 381454
rect 452382 380898 452414 381454
rect 451794 345454 452414 380898
rect 451794 344898 451826 345454
rect 452382 344898 452414 345454
rect 451794 309454 452414 344898
rect 451794 308898 451826 309454
rect 452382 308898 452414 309454
rect 451794 273454 452414 308898
rect 451794 272898 451826 273454
rect 452382 272898 452414 273454
rect 451794 237454 452414 272898
rect 451794 236898 451826 237454
rect 452382 236898 452414 237454
rect 451794 201454 452414 236898
rect 451794 200898 451826 201454
rect 452382 200898 452414 201454
rect 451794 165454 452414 200898
rect 451794 164898 451826 165454
rect 452382 164898 452414 165454
rect 451794 129454 452414 164898
rect 451794 128898 451826 129454
rect 452382 128898 452414 129454
rect 451794 93454 452414 128898
rect 451794 92898 451826 93454
rect 452382 92898 452414 93454
rect 451794 57454 452414 92898
rect 451794 56898 451826 57454
rect 452382 56898 452414 57454
rect 451794 21454 452414 56898
rect 451794 20898 451826 21454
rect 452382 20898 452414 21454
rect 451794 -1306 452414 20898
rect 451794 -1862 451826 -1306
rect 452382 -1862 452414 -1306
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672618 455546 673174
rect 456102 672618 456134 673174
rect 455514 637174 456134 672618
rect 455514 636618 455546 637174
rect 456102 636618 456134 637174
rect 455514 601174 456134 636618
rect 455514 600618 455546 601174
rect 456102 600618 456134 601174
rect 455514 565174 456134 600618
rect 455514 564618 455546 565174
rect 456102 564618 456134 565174
rect 455514 529174 456134 564618
rect 455514 528618 455546 529174
rect 456102 528618 456134 529174
rect 455514 493174 456134 528618
rect 455514 492618 455546 493174
rect 456102 492618 456134 493174
rect 455514 457174 456134 492618
rect 455514 456618 455546 457174
rect 456102 456618 456134 457174
rect 455514 421174 456134 456618
rect 455514 420618 455546 421174
rect 456102 420618 456134 421174
rect 455514 385174 456134 420618
rect 455514 384618 455546 385174
rect 456102 384618 456134 385174
rect 455514 349174 456134 384618
rect 455514 348618 455546 349174
rect 456102 348618 456134 349174
rect 455514 313174 456134 348618
rect 455514 312618 455546 313174
rect 456102 312618 456134 313174
rect 455514 277174 456134 312618
rect 455514 276618 455546 277174
rect 456102 276618 456134 277174
rect 455514 241174 456134 276618
rect 455514 240618 455546 241174
rect 456102 240618 456134 241174
rect 455514 205174 456134 240618
rect 455514 204618 455546 205174
rect 456102 204618 456134 205174
rect 455514 169174 456134 204618
rect 455514 168618 455546 169174
rect 456102 168618 456134 169174
rect 455514 133174 456134 168618
rect 455514 132618 455546 133174
rect 456102 132618 456134 133174
rect 455514 97174 456134 132618
rect 455514 96618 455546 97174
rect 456102 96618 456134 97174
rect 455514 61174 456134 96618
rect 455514 60618 455546 61174
rect 456102 60618 456134 61174
rect 455514 25174 456134 60618
rect 455514 24618 455546 25174
rect 456102 24618 456134 25174
rect 455514 -3226 456134 24618
rect 455514 -3782 455546 -3226
rect 456102 -3782 456134 -3226
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676338 459266 676894
rect 459822 676338 459854 676894
rect 459234 640894 459854 676338
rect 459234 640338 459266 640894
rect 459822 640338 459854 640894
rect 459234 604894 459854 640338
rect 459234 604338 459266 604894
rect 459822 604338 459854 604894
rect 459234 568894 459854 604338
rect 459234 568338 459266 568894
rect 459822 568338 459854 568894
rect 459234 532894 459854 568338
rect 459234 532338 459266 532894
rect 459822 532338 459854 532894
rect 459234 496894 459854 532338
rect 459234 496338 459266 496894
rect 459822 496338 459854 496894
rect 459234 460894 459854 496338
rect 459234 460338 459266 460894
rect 459822 460338 459854 460894
rect 459234 424894 459854 460338
rect 459234 424338 459266 424894
rect 459822 424338 459854 424894
rect 459234 388894 459854 424338
rect 459234 388338 459266 388894
rect 459822 388338 459854 388894
rect 459234 352894 459854 388338
rect 459234 352338 459266 352894
rect 459822 352338 459854 352894
rect 459234 316894 459854 352338
rect 459234 316338 459266 316894
rect 459822 316338 459854 316894
rect 459234 280894 459854 316338
rect 459234 280338 459266 280894
rect 459822 280338 459854 280894
rect 459234 244894 459854 280338
rect 459234 244338 459266 244894
rect 459822 244338 459854 244894
rect 459234 208894 459854 244338
rect 459234 208338 459266 208894
rect 459822 208338 459854 208894
rect 459234 172894 459854 208338
rect 459234 172338 459266 172894
rect 459822 172338 459854 172894
rect 459234 136894 459854 172338
rect 459234 136338 459266 136894
rect 459822 136338 459854 136894
rect 459234 100894 459854 136338
rect 459234 100338 459266 100894
rect 459822 100338 459854 100894
rect 459234 64894 459854 100338
rect 459234 64338 459266 64894
rect 459822 64338 459854 64894
rect 459234 28894 459854 64338
rect 459234 28338 459266 28894
rect 459822 28338 459854 28894
rect 459234 -5146 459854 28338
rect 459234 -5702 459266 -5146
rect 459822 -5702 459854 -5146
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710042 480986 710598
rect 481542 710042 481574 710598
rect 477234 708678 477854 709670
rect 477234 708122 477266 708678
rect 477822 708122 477854 708678
rect 473514 706758 474134 707750
rect 473514 706202 473546 706758
rect 474102 706202 474134 706758
rect 462954 680058 462986 680614
rect 463542 680058 463574 680614
rect 462954 644614 463574 680058
rect 462954 644058 462986 644614
rect 463542 644058 463574 644614
rect 462954 608614 463574 644058
rect 462954 608058 462986 608614
rect 463542 608058 463574 608614
rect 462954 572614 463574 608058
rect 462954 572058 462986 572614
rect 463542 572058 463574 572614
rect 462954 536614 463574 572058
rect 462954 536058 462986 536614
rect 463542 536058 463574 536614
rect 462954 500614 463574 536058
rect 462954 500058 462986 500614
rect 463542 500058 463574 500614
rect 462954 464614 463574 500058
rect 462954 464058 462986 464614
rect 463542 464058 463574 464614
rect 462954 428614 463574 464058
rect 462954 428058 462986 428614
rect 463542 428058 463574 428614
rect 462954 392614 463574 428058
rect 462954 392058 462986 392614
rect 463542 392058 463574 392614
rect 462954 356614 463574 392058
rect 462954 356058 462986 356614
rect 463542 356058 463574 356614
rect 462954 320614 463574 356058
rect 462954 320058 462986 320614
rect 463542 320058 463574 320614
rect 462954 284614 463574 320058
rect 462954 284058 462986 284614
rect 463542 284058 463574 284614
rect 462954 248614 463574 284058
rect 462954 248058 462986 248614
rect 463542 248058 463574 248614
rect 462954 212614 463574 248058
rect 462954 212058 462986 212614
rect 463542 212058 463574 212614
rect 462954 176614 463574 212058
rect 462954 176058 462986 176614
rect 463542 176058 463574 176614
rect 462954 140614 463574 176058
rect 462954 140058 462986 140614
rect 463542 140058 463574 140614
rect 462954 104614 463574 140058
rect 462954 104058 462986 104614
rect 463542 104058 463574 104614
rect 462954 68614 463574 104058
rect 462954 68058 462986 68614
rect 463542 68058 463574 68614
rect 462954 32614 463574 68058
rect 462954 32058 462986 32614
rect 463542 32058 463574 32614
rect 444954 -6662 444986 -6106
rect 445542 -6662 445574 -6106
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704282 469826 704838
rect 470382 704282 470414 704838
rect 469794 687454 470414 704282
rect 469794 686898 469826 687454
rect 470382 686898 470414 687454
rect 469794 651454 470414 686898
rect 469794 650898 469826 651454
rect 470382 650898 470414 651454
rect 469794 615454 470414 650898
rect 469794 614898 469826 615454
rect 470382 614898 470414 615454
rect 469794 579454 470414 614898
rect 469794 578898 469826 579454
rect 470382 578898 470414 579454
rect 469794 543454 470414 578898
rect 469794 542898 469826 543454
rect 470382 542898 470414 543454
rect 469794 507454 470414 542898
rect 469794 506898 469826 507454
rect 470382 506898 470414 507454
rect 469794 471454 470414 506898
rect 469794 470898 469826 471454
rect 470382 470898 470414 471454
rect 469794 435454 470414 470898
rect 469794 434898 469826 435454
rect 470382 434898 470414 435454
rect 469794 399454 470414 434898
rect 469794 398898 469826 399454
rect 470382 398898 470414 399454
rect 469794 363454 470414 398898
rect 469794 362898 469826 363454
rect 470382 362898 470414 363454
rect 469794 327454 470414 362898
rect 469794 326898 469826 327454
rect 470382 326898 470414 327454
rect 469794 291454 470414 326898
rect 469794 290898 469826 291454
rect 470382 290898 470414 291454
rect 469794 255454 470414 290898
rect 469794 254898 469826 255454
rect 470382 254898 470414 255454
rect 469794 219454 470414 254898
rect 469794 218898 469826 219454
rect 470382 218898 470414 219454
rect 469794 183454 470414 218898
rect 469794 182898 469826 183454
rect 470382 182898 470414 183454
rect 469794 147454 470414 182898
rect 469794 146898 469826 147454
rect 470382 146898 470414 147454
rect 469794 111454 470414 146898
rect 469794 110898 469826 111454
rect 470382 110898 470414 111454
rect 469794 75454 470414 110898
rect 469794 74898 469826 75454
rect 470382 74898 470414 75454
rect 469794 39454 470414 74898
rect 469794 38898 469826 39454
rect 470382 38898 470414 39454
rect 469794 3454 470414 38898
rect 469794 2898 469826 3454
rect 470382 2898 470414 3454
rect 469794 -346 470414 2898
rect 469794 -902 469826 -346
rect 470382 -902 470414 -346
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690618 473546 691174
rect 474102 690618 474134 691174
rect 473514 655174 474134 690618
rect 473514 654618 473546 655174
rect 474102 654618 474134 655174
rect 473514 619174 474134 654618
rect 473514 618618 473546 619174
rect 474102 618618 474134 619174
rect 473514 583174 474134 618618
rect 473514 582618 473546 583174
rect 474102 582618 474134 583174
rect 473514 547174 474134 582618
rect 473514 546618 473546 547174
rect 474102 546618 474134 547174
rect 473514 511174 474134 546618
rect 473514 510618 473546 511174
rect 474102 510618 474134 511174
rect 473514 475174 474134 510618
rect 473514 474618 473546 475174
rect 474102 474618 474134 475174
rect 473514 439174 474134 474618
rect 473514 438618 473546 439174
rect 474102 438618 474134 439174
rect 473514 403174 474134 438618
rect 473514 402618 473546 403174
rect 474102 402618 474134 403174
rect 473514 367174 474134 402618
rect 473514 366618 473546 367174
rect 474102 366618 474134 367174
rect 473514 331174 474134 366618
rect 473514 330618 473546 331174
rect 474102 330618 474134 331174
rect 473514 295174 474134 330618
rect 473514 294618 473546 295174
rect 474102 294618 474134 295174
rect 473514 259174 474134 294618
rect 473514 258618 473546 259174
rect 474102 258618 474134 259174
rect 473514 223174 474134 258618
rect 473514 222618 473546 223174
rect 474102 222618 474134 223174
rect 473514 187174 474134 222618
rect 473514 186618 473546 187174
rect 474102 186618 474134 187174
rect 473514 151174 474134 186618
rect 473514 150618 473546 151174
rect 474102 150618 474134 151174
rect 473514 115174 474134 150618
rect 473514 114618 473546 115174
rect 474102 114618 474134 115174
rect 473514 79174 474134 114618
rect 473514 78618 473546 79174
rect 474102 78618 474134 79174
rect 473514 43174 474134 78618
rect 473514 42618 473546 43174
rect 474102 42618 474134 43174
rect 473514 7174 474134 42618
rect 473514 6618 473546 7174
rect 474102 6618 474134 7174
rect 473514 -2266 474134 6618
rect 473514 -2822 473546 -2266
rect 474102 -2822 474134 -2266
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694338 477266 694894
rect 477822 694338 477854 694894
rect 477234 658894 477854 694338
rect 477234 658338 477266 658894
rect 477822 658338 477854 658894
rect 477234 622894 477854 658338
rect 477234 622338 477266 622894
rect 477822 622338 477854 622894
rect 477234 586894 477854 622338
rect 477234 586338 477266 586894
rect 477822 586338 477854 586894
rect 477234 550894 477854 586338
rect 477234 550338 477266 550894
rect 477822 550338 477854 550894
rect 477234 514894 477854 550338
rect 477234 514338 477266 514894
rect 477822 514338 477854 514894
rect 477234 478894 477854 514338
rect 477234 478338 477266 478894
rect 477822 478338 477854 478894
rect 477234 442894 477854 478338
rect 477234 442338 477266 442894
rect 477822 442338 477854 442894
rect 477234 406894 477854 442338
rect 477234 406338 477266 406894
rect 477822 406338 477854 406894
rect 477234 370894 477854 406338
rect 477234 370338 477266 370894
rect 477822 370338 477854 370894
rect 477234 334894 477854 370338
rect 477234 334338 477266 334894
rect 477822 334338 477854 334894
rect 477234 298894 477854 334338
rect 477234 298338 477266 298894
rect 477822 298338 477854 298894
rect 477234 262894 477854 298338
rect 477234 262338 477266 262894
rect 477822 262338 477854 262894
rect 477234 226894 477854 262338
rect 477234 226338 477266 226894
rect 477822 226338 477854 226894
rect 477234 190894 477854 226338
rect 477234 190338 477266 190894
rect 477822 190338 477854 190894
rect 477234 154894 477854 190338
rect 477234 154338 477266 154894
rect 477822 154338 477854 154894
rect 477234 118894 477854 154338
rect 477234 118338 477266 118894
rect 477822 118338 477854 118894
rect 477234 82894 477854 118338
rect 477234 82338 477266 82894
rect 477822 82338 477854 82894
rect 477234 46894 477854 82338
rect 477234 46338 477266 46894
rect 477822 46338 477854 46894
rect 477234 10894 477854 46338
rect 477234 10338 477266 10894
rect 477822 10338 477854 10894
rect 477234 -4186 477854 10338
rect 477234 -4742 477266 -4186
rect 477822 -4742 477854 -4186
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711002 498986 711558
rect 499542 711002 499574 711558
rect 495234 709638 495854 709670
rect 495234 709082 495266 709638
rect 495822 709082 495854 709638
rect 491514 707718 492134 707750
rect 491514 707162 491546 707718
rect 492102 707162 492134 707718
rect 480954 698058 480986 698614
rect 481542 698058 481574 698614
rect 480954 662614 481574 698058
rect 480954 662058 480986 662614
rect 481542 662058 481574 662614
rect 480954 626614 481574 662058
rect 480954 626058 480986 626614
rect 481542 626058 481574 626614
rect 480954 590614 481574 626058
rect 480954 590058 480986 590614
rect 481542 590058 481574 590614
rect 480954 554614 481574 590058
rect 480954 554058 480986 554614
rect 481542 554058 481574 554614
rect 480954 518614 481574 554058
rect 480954 518058 480986 518614
rect 481542 518058 481574 518614
rect 480954 482614 481574 518058
rect 480954 482058 480986 482614
rect 481542 482058 481574 482614
rect 480954 446614 481574 482058
rect 480954 446058 480986 446614
rect 481542 446058 481574 446614
rect 480954 410614 481574 446058
rect 480954 410058 480986 410614
rect 481542 410058 481574 410614
rect 480954 374614 481574 410058
rect 480954 374058 480986 374614
rect 481542 374058 481574 374614
rect 480954 338614 481574 374058
rect 480954 338058 480986 338614
rect 481542 338058 481574 338614
rect 480954 302614 481574 338058
rect 480954 302058 480986 302614
rect 481542 302058 481574 302614
rect 480954 266614 481574 302058
rect 480954 266058 480986 266614
rect 481542 266058 481574 266614
rect 480954 230614 481574 266058
rect 480954 230058 480986 230614
rect 481542 230058 481574 230614
rect 480954 194614 481574 230058
rect 480954 194058 480986 194614
rect 481542 194058 481574 194614
rect 480954 158614 481574 194058
rect 480954 158058 480986 158614
rect 481542 158058 481574 158614
rect 480954 122614 481574 158058
rect 480954 122058 480986 122614
rect 481542 122058 481574 122614
rect 480954 86614 481574 122058
rect 480954 86058 480986 86614
rect 481542 86058 481574 86614
rect 480954 50614 481574 86058
rect 480954 50058 480986 50614
rect 481542 50058 481574 50614
rect 480954 14614 481574 50058
rect 480954 14058 480986 14614
rect 481542 14058 481574 14614
rect 462954 -7622 462986 -7066
rect 463542 -7622 463574 -7066
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705242 487826 705798
rect 488382 705242 488414 705798
rect 487794 669454 488414 705242
rect 487794 668898 487826 669454
rect 488382 668898 488414 669454
rect 487794 633454 488414 668898
rect 487794 632898 487826 633454
rect 488382 632898 488414 633454
rect 487794 597454 488414 632898
rect 487794 596898 487826 597454
rect 488382 596898 488414 597454
rect 487794 561454 488414 596898
rect 487794 560898 487826 561454
rect 488382 560898 488414 561454
rect 487794 525454 488414 560898
rect 487794 524898 487826 525454
rect 488382 524898 488414 525454
rect 487794 489454 488414 524898
rect 487794 488898 487826 489454
rect 488382 488898 488414 489454
rect 487794 453454 488414 488898
rect 487794 452898 487826 453454
rect 488382 452898 488414 453454
rect 487794 417454 488414 452898
rect 487794 416898 487826 417454
rect 488382 416898 488414 417454
rect 487794 381454 488414 416898
rect 487794 380898 487826 381454
rect 488382 380898 488414 381454
rect 487794 345454 488414 380898
rect 487794 344898 487826 345454
rect 488382 344898 488414 345454
rect 487794 309454 488414 344898
rect 487794 308898 487826 309454
rect 488382 308898 488414 309454
rect 487794 273454 488414 308898
rect 487794 272898 487826 273454
rect 488382 272898 488414 273454
rect 487794 237454 488414 272898
rect 487794 236898 487826 237454
rect 488382 236898 488414 237454
rect 487794 201454 488414 236898
rect 487794 200898 487826 201454
rect 488382 200898 488414 201454
rect 487794 165454 488414 200898
rect 487794 164898 487826 165454
rect 488382 164898 488414 165454
rect 487794 129454 488414 164898
rect 487794 128898 487826 129454
rect 488382 128898 488414 129454
rect 487794 93454 488414 128898
rect 487794 92898 487826 93454
rect 488382 92898 488414 93454
rect 487794 57454 488414 92898
rect 487794 56898 487826 57454
rect 488382 56898 488414 57454
rect 487794 21454 488414 56898
rect 487794 20898 487826 21454
rect 488382 20898 488414 21454
rect 487794 -1306 488414 20898
rect 487794 -1862 487826 -1306
rect 488382 -1862 488414 -1306
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672618 491546 673174
rect 492102 672618 492134 673174
rect 491514 637174 492134 672618
rect 491514 636618 491546 637174
rect 492102 636618 492134 637174
rect 491514 601174 492134 636618
rect 491514 600618 491546 601174
rect 492102 600618 492134 601174
rect 491514 565174 492134 600618
rect 491514 564618 491546 565174
rect 492102 564618 492134 565174
rect 491514 529174 492134 564618
rect 491514 528618 491546 529174
rect 492102 528618 492134 529174
rect 491514 493174 492134 528618
rect 491514 492618 491546 493174
rect 492102 492618 492134 493174
rect 491514 457174 492134 492618
rect 491514 456618 491546 457174
rect 492102 456618 492134 457174
rect 491514 421174 492134 456618
rect 491514 420618 491546 421174
rect 492102 420618 492134 421174
rect 491514 385174 492134 420618
rect 491514 384618 491546 385174
rect 492102 384618 492134 385174
rect 491514 349174 492134 384618
rect 491514 348618 491546 349174
rect 492102 348618 492134 349174
rect 491514 313174 492134 348618
rect 491514 312618 491546 313174
rect 492102 312618 492134 313174
rect 491514 277174 492134 312618
rect 491514 276618 491546 277174
rect 492102 276618 492134 277174
rect 491514 241174 492134 276618
rect 491514 240618 491546 241174
rect 492102 240618 492134 241174
rect 491514 205174 492134 240618
rect 491514 204618 491546 205174
rect 492102 204618 492134 205174
rect 491514 169174 492134 204618
rect 491514 168618 491546 169174
rect 492102 168618 492134 169174
rect 491514 133174 492134 168618
rect 491514 132618 491546 133174
rect 492102 132618 492134 133174
rect 491514 97174 492134 132618
rect 491514 96618 491546 97174
rect 492102 96618 492134 97174
rect 491514 61174 492134 96618
rect 491514 60618 491546 61174
rect 492102 60618 492134 61174
rect 491514 25174 492134 60618
rect 491514 24618 491546 25174
rect 492102 24618 492134 25174
rect 491514 -3226 492134 24618
rect 491514 -3782 491546 -3226
rect 492102 -3782 492134 -3226
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676338 495266 676894
rect 495822 676338 495854 676894
rect 495234 640894 495854 676338
rect 495234 640338 495266 640894
rect 495822 640338 495854 640894
rect 495234 604894 495854 640338
rect 495234 604338 495266 604894
rect 495822 604338 495854 604894
rect 495234 568894 495854 604338
rect 495234 568338 495266 568894
rect 495822 568338 495854 568894
rect 495234 532894 495854 568338
rect 495234 532338 495266 532894
rect 495822 532338 495854 532894
rect 495234 496894 495854 532338
rect 495234 496338 495266 496894
rect 495822 496338 495854 496894
rect 495234 460894 495854 496338
rect 495234 460338 495266 460894
rect 495822 460338 495854 460894
rect 495234 424894 495854 460338
rect 495234 424338 495266 424894
rect 495822 424338 495854 424894
rect 495234 388894 495854 424338
rect 495234 388338 495266 388894
rect 495822 388338 495854 388894
rect 495234 352894 495854 388338
rect 495234 352338 495266 352894
rect 495822 352338 495854 352894
rect 495234 316894 495854 352338
rect 495234 316338 495266 316894
rect 495822 316338 495854 316894
rect 495234 280894 495854 316338
rect 495234 280338 495266 280894
rect 495822 280338 495854 280894
rect 495234 244894 495854 280338
rect 495234 244338 495266 244894
rect 495822 244338 495854 244894
rect 495234 208894 495854 244338
rect 495234 208338 495266 208894
rect 495822 208338 495854 208894
rect 495234 172894 495854 208338
rect 495234 172338 495266 172894
rect 495822 172338 495854 172894
rect 495234 136894 495854 172338
rect 495234 136338 495266 136894
rect 495822 136338 495854 136894
rect 495234 100894 495854 136338
rect 495234 100338 495266 100894
rect 495822 100338 495854 100894
rect 495234 64894 495854 100338
rect 495234 64338 495266 64894
rect 495822 64338 495854 64894
rect 495234 28894 495854 64338
rect 495234 28338 495266 28894
rect 495822 28338 495854 28894
rect 495234 -5146 495854 28338
rect 495234 -5702 495266 -5146
rect 495822 -5702 495854 -5146
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710042 516986 710598
rect 517542 710042 517574 710598
rect 513234 708678 513854 709670
rect 513234 708122 513266 708678
rect 513822 708122 513854 708678
rect 509514 706758 510134 707750
rect 509514 706202 509546 706758
rect 510102 706202 510134 706758
rect 498954 680058 498986 680614
rect 499542 680058 499574 680614
rect 498954 644614 499574 680058
rect 498954 644058 498986 644614
rect 499542 644058 499574 644614
rect 498954 608614 499574 644058
rect 498954 608058 498986 608614
rect 499542 608058 499574 608614
rect 498954 572614 499574 608058
rect 498954 572058 498986 572614
rect 499542 572058 499574 572614
rect 498954 536614 499574 572058
rect 498954 536058 498986 536614
rect 499542 536058 499574 536614
rect 498954 500614 499574 536058
rect 498954 500058 498986 500614
rect 499542 500058 499574 500614
rect 498954 464614 499574 500058
rect 498954 464058 498986 464614
rect 499542 464058 499574 464614
rect 498954 428614 499574 464058
rect 498954 428058 498986 428614
rect 499542 428058 499574 428614
rect 498954 392614 499574 428058
rect 498954 392058 498986 392614
rect 499542 392058 499574 392614
rect 498954 356614 499574 392058
rect 498954 356058 498986 356614
rect 499542 356058 499574 356614
rect 498954 320614 499574 356058
rect 498954 320058 498986 320614
rect 499542 320058 499574 320614
rect 498954 284614 499574 320058
rect 498954 284058 498986 284614
rect 499542 284058 499574 284614
rect 498954 248614 499574 284058
rect 498954 248058 498986 248614
rect 499542 248058 499574 248614
rect 498954 212614 499574 248058
rect 498954 212058 498986 212614
rect 499542 212058 499574 212614
rect 498954 176614 499574 212058
rect 498954 176058 498986 176614
rect 499542 176058 499574 176614
rect 498954 140614 499574 176058
rect 498954 140058 498986 140614
rect 499542 140058 499574 140614
rect 498954 104614 499574 140058
rect 498954 104058 498986 104614
rect 499542 104058 499574 104614
rect 498954 68614 499574 104058
rect 498954 68058 498986 68614
rect 499542 68058 499574 68614
rect 498954 32614 499574 68058
rect 498954 32058 498986 32614
rect 499542 32058 499574 32614
rect 480954 -6662 480986 -6106
rect 481542 -6662 481574 -6106
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704282 505826 704838
rect 506382 704282 506414 704838
rect 505794 687454 506414 704282
rect 505794 686898 505826 687454
rect 506382 686898 506414 687454
rect 505794 651454 506414 686898
rect 505794 650898 505826 651454
rect 506382 650898 506414 651454
rect 505794 615454 506414 650898
rect 505794 614898 505826 615454
rect 506382 614898 506414 615454
rect 505794 579454 506414 614898
rect 505794 578898 505826 579454
rect 506382 578898 506414 579454
rect 505794 543454 506414 578898
rect 505794 542898 505826 543454
rect 506382 542898 506414 543454
rect 505794 507454 506414 542898
rect 505794 506898 505826 507454
rect 506382 506898 506414 507454
rect 505794 471454 506414 506898
rect 505794 470898 505826 471454
rect 506382 470898 506414 471454
rect 505794 435454 506414 470898
rect 505794 434898 505826 435454
rect 506382 434898 506414 435454
rect 505794 399454 506414 434898
rect 505794 398898 505826 399454
rect 506382 398898 506414 399454
rect 505794 363454 506414 398898
rect 505794 362898 505826 363454
rect 506382 362898 506414 363454
rect 505794 327454 506414 362898
rect 505794 326898 505826 327454
rect 506382 326898 506414 327454
rect 505794 291454 506414 326898
rect 505794 290898 505826 291454
rect 506382 290898 506414 291454
rect 505794 255454 506414 290898
rect 505794 254898 505826 255454
rect 506382 254898 506414 255454
rect 505794 219454 506414 254898
rect 505794 218898 505826 219454
rect 506382 218898 506414 219454
rect 505794 183454 506414 218898
rect 505794 182898 505826 183454
rect 506382 182898 506414 183454
rect 505794 147454 506414 182898
rect 505794 146898 505826 147454
rect 506382 146898 506414 147454
rect 505794 111454 506414 146898
rect 505794 110898 505826 111454
rect 506382 110898 506414 111454
rect 505794 75454 506414 110898
rect 505794 74898 505826 75454
rect 506382 74898 506414 75454
rect 505794 39454 506414 74898
rect 505794 38898 505826 39454
rect 506382 38898 506414 39454
rect 505794 3454 506414 38898
rect 505794 2898 505826 3454
rect 506382 2898 506414 3454
rect 505794 -346 506414 2898
rect 505794 -902 505826 -346
rect 506382 -902 506414 -346
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690618 509546 691174
rect 510102 690618 510134 691174
rect 509514 655174 510134 690618
rect 509514 654618 509546 655174
rect 510102 654618 510134 655174
rect 509514 619174 510134 654618
rect 509514 618618 509546 619174
rect 510102 618618 510134 619174
rect 509514 583174 510134 618618
rect 509514 582618 509546 583174
rect 510102 582618 510134 583174
rect 509514 547174 510134 582618
rect 509514 546618 509546 547174
rect 510102 546618 510134 547174
rect 509514 511174 510134 546618
rect 509514 510618 509546 511174
rect 510102 510618 510134 511174
rect 509514 475174 510134 510618
rect 509514 474618 509546 475174
rect 510102 474618 510134 475174
rect 509514 439174 510134 474618
rect 509514 438618 509546 439174
rect 510102 438618 510134 439174
rect 509514 403174 510134 438618
rect 509514 402618 509546 403174
rect 510102 402618 510134 403174
rect 509514 367174 510134 402618
rect 509514 366618 509546 367174
rect 510102 366618 510134 367174
rect 509514 331174 510134 366618
rect 509514 330618 509546 331174
rect 510102 330618 510134 331174
rect 509514 295174 510134 330618
rect 509514 294618 509546 295174
rect 510102 294618 510134 295174
rect 509514 259174 510134 294618
rect 509514 258618 509546 259174
rect 510102 258618 510134 259174
rect 509514 223174 510134 258618
rect 509514 222618 509546 223174
rect 510102 222618 510134 223174
rect 509514 187174 510134 222618
rect 509514 186618 509546 187174
rect 510102 186618 510134 187174
rect 509514 151174 510134 186618
rect 509514 150618 509546 151174
rect 510102 150618 510134 151174
rect 509514 115174 510134 150618
rect 509514 114618 509546 115174
rect 510102 114618 510134 115174
rect 509514 79174 510134 114618
rect 509514 78618 509546 79174
rect 510102 78618 510134 79174
rect 509514 43174 510134 78618
rect 509514 42618 509546 43174
rect 510102 42618 510134 43174
rect 509514 7174 510134 42618
rect 509514 6618 509546 7174
rect 510102 6618 510134 7174
rect 509514 -2266 510134 6618
rect 509514 -2822 509546 -2266
rect 510102 -2822 510134 -2266
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694338 513266 694894
rect 513822 694338 513854 694894
rect 513234 658894 513854 694338
rect 513234 658338 513266 658894
rect 513822 658338 513854 658894
rect 513234 622894 513854 658338
rect 513234 622338 513266 622894
rect 513822 622338 513854 622894
rect 513234 586894 513854 622338
rect 513234 586338 513266 586894
rect 513822 586338 513854 586894
rect 513234 550894 513854 586338
rect 513234 550338 513266 550894
rect 513822 550338 513854 550894
rect 513234 514894 513854 550338
rect 513234 514338 513266 514894
rect 513822 514338 513854 514894
rect 513234 478894 513854 514338
rect 513234 478338 513266 478894
rect 513822 478338 513854 478894
rect 513234 442894 513854 478338
rect 513234 442338 513266 442894
rect 513822 442338 513854 442894
rect 513234 406894 513854 442338
rect 513234 406338 513266 406894
rect 513822 406338 513854 406894
rect 513234 370894 513854 406338
rect 513234 370338 513266 370894
rect 513822 370338 513854 370894
rect 513234 334894 513854 370338
rect 513234 334338 513266 334894
rect 513822 334338 513854 334894
rect 513234 298894 513854 334338
rect 513234 298338 513266 298894
rect 513822 298338 513854 298894
rect 513234 262894 513854 298338
rect 513234 262338 513266 262894
rect 513822 262338 513854 262894
rect 513234 226894 513854 262338
rect 513234 226338 513266 226894
rect 513822 226338 513854 226894
rect 513234 190894 513854 226338
rect 513234 190338 513266 190894
rect 513822 190338 513854 190894
rect 513234 154894 513854 190338
rect 513234 154338 513266 154894
rect 513822 154338 513854 154894
rect 513234 118894 513854 154338
rect 513234 118338 513266 118894
rect 513822 118338 513854 118894
rect 513234 82894 513854 118338
rect 513234 82338 513266 82894
rect 513822 82338 513854 82894
rect 513234 46894 513854 82338
rect 513234 46338 513266 46894
rect 513822 46338 513854 46894
rect 513234 10894 513854 46338
rect 513234 10338 513266 10894
rect 513822 10338 513854 10894
rect 513234 -4186 513854 10338
rect 513234 -4742 513266 -4186
rect 513822 -4742 513854 -4186
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711002 534986 711558
rect 535542 711002 535574 711558
rect 531234 709638 531854 709670
rect 531234 709082 531266 709638
rect 531822 709082 531854 709638
rect 527514 707718 528134 707750
rect 527514 707162 527546 707718
rect 528102 707162 528134 707718
rect 516954 698058 516986 698614
rect 517542 698058 517574 698614
rect 516954 662614 517574 698058
rect 516954 662058 516986 662614
rect 517542 662058 517574 662614
rect 516954 626614 517574 662058
rect 516954 626058 516986 626614
rect 517542 626058 517574 626614
rect 516954 590614 517574 626058
rect 516954 590058 516986 590614
rect 517542 590058 517574 590614
rect 516954 554614 517574 590058
rect 516954 554058 516986 554614
rect 517542 554058 517574 554614
rect 516954 518614 517574 554058
rect 516954 518058 516986 518614
rect 517542 518058 517574 518614
rect 516954 482614 517574 518058
rect 516954 482058 516986 482614
rect 517542 482058 517574 482614
rect 516954 446614 517574 482058
rect 516954 446058 516986 446614
rect 517542 446058 517574 446614
rect 516954 410614 517574 446058
rect 516954 410058 516986 410614
rect 517542 410058 517574 410614
rect 516954 374614 517574 410058
rect 516954 374058 516986 374614
rect 517542 374058 517574 374614
rect 516954 338614 517574 374058
rect 516954 338058 516986 338614
rect 517542 338058 517574 338614
rect 516954 302614 517574 338058
rect 516954 302058 516986 302614
rect 517542 302058 517574 302614
rect 516954 266614 517574 302058
rect 516954 266058 516986 266614
rect 517542 266058 517574 266614
rect 516954 230614 517574 266058
rect 516954 230058 516986 230614
rect 517542 230058 517574 230614
rect 516954 194614 517574 230058
rect 516954 194058 516986 194614
rect 517542 194058 517574 194614
rect 516954 158614 517574 194058
rect 516954 158058 516986 158614
rect 517542 158058 517574 158614
rect 516954 122614 517574 158058
rect 516954 122058 516986 122614
rect 517542 122058 517574 122614
rect 516954 86614 517574 122058
rect 516954 86058 516986 86614
rect 517542 86058 517574 86614
rect 516954 50614 517574 86058
rect 516954 50058 516986 50614
rect 517542 50058 517574 50614
rect 516954 14614 517574 50058
rect 516954 14058 516986 14614
rect 517542 14058 517574 14614
rect 498954 -7622 498986 -7066
rect 499542 -7622 499574 -7066
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705242 523826 705798
rect 524382 705242 524414 705798
rect 523794 669454 524414 705242
rect 523794 668898 523826 669454
rect 524382 668898 524414 669454
rect 523794 633454 524414 668898
rect 523794 632898 523826 633454
rect 524382 632898 524414 633454
rect 523794 597454 524414 632898
rect 523794 596898 523826 597454
rect 524382 596898 524414 597454
rect 523794 561454 524414 596898
rect 523794 560898 523826 561454
rect 524382 560898 524414 561454
rect 523794 525454 524414 560898
rect 523794 524898 523826 525454
rect 524382 524898 524414 525454
rect 523794 489454 524414 524898
rect 523794 488898 523826 489454
rect 524382 488898 524414 489454
rect 523794 453454 524414 488898
rect 523794 452898 523826 453454
rect 524382 452898 524414 453454
rect 523794 417454 524414 452898
rect 523794 416898 523826 417454
rect 524382 416898 524414 417454
rect 523794 381454 524414 416898
rect 523794 380898 523826 381454
rect 524382 380898 524414 381454
rect 523794 345454 524414 380898
rect 523794 344898 523826 345454
rect 524382 344898 524414 345454
rect 523794 309454 524414 344898
rect 523794 308898 523826 309454
rect 524382 308898 524414 309454
rect 523794 273454 524414 308898
rect 523794 272898 523826 273454
rect 524382 272898 524414 273454
rect 523794 237454 524414 272898
rect 523794 236898 523826 237454
rect 524382 236898 524414 237454
rect 523794 201454 524414 236898
rect 523794 200898 523826 201454
rect 524382 200898 524414 201454
rect 523794 165454 524414 200898
rect 523794 164898 523826 165454
rect 524382 164898 524414 165454
rect 523794 129454 524414 164898
rect 523794 128898 523826 129454
rect 524382 128898 524414 129454
rect 523794 93454 524414 128898
rect 523794 92898 523826 93454
rect 524382 92898 524414 93454
rect 523794 57454 524414 92898
rect 523794 56898 523826 57454
rect 524382 56898 524414 57454
rect 523794 21454 524414 56898
rect 523794 20898 523826 21454
rect 524382 20898 524414 21454
rect 523794 -1306 524414 20898
rect 523794 -1862 523826 -1306
rect 524382 -1862 524414 -1306
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672618 527546 673174
rect 528102 672618 528134 673174
rect 527514 637174 528134 672618
rect 527514 636618 527546 637174
rect 528102 636618 528134 637174
rect 527514 601174 528134 636618
rect 527514 600618 527546 601174
rect 528102 600618 528134 601174
rect 527514 565174 528134 600618
rect 527514 564618 527546 565174
rect 528102 564618 528134 565174
rect 527514 529174 528134 564618
rect 527514 528618 527546 529174
rect 528102 528618 528134 529174
rect 527514 493174 528134 528618
rect 527514 492618 527546 493174
rect 528102 492618 528134 493174
rect 527514 457174 528134 492618
rect 527514 456618 527546 457174
rect 528102 456618 528134 457174
rect 527514 421174 528134 456618
rect 527514 420618 527546 421174
rect 528102 420618 528134 421174
rect 527514 385174 528134 420618
rect 527514 384618 527546 385174
rect 528102 384618 528134 385174
rect 527514 349174 528134 384618
rect 527514 348618 527546 349174
rect 528102 348618 528134 349174
rect 527514 313174 528134 348618
rect 527514 312618 527546 313174
rect 528102 312618 528134 313174
rect 527514 277174 528134 312618
rect 527514 276618 527546 277174
rect 528102 276618 528134 277174
rect 527514 241174 528134 276618
rect 527514 240618 527546 241174
rect 528102 240618 528134 241174
rect 527514 205174 528134 240618
rect 527514 204618 527546 205174
rect 528102 204618 528134 205174
rect 527514 169174 528134 204618
rect 527514 168618 527546 169174
rect 528102 168618 528134 169174
rect 527514 133174 528134 168618
rect 527514 132618 527546 133174
rect 528102 132618 528134 133174
rect 527514 97174 528134 132618
rect 527514 96618 527546 97174
rect 528102 96618 528134 97174
rect 527514 61174 528134 96618
rect 527514 60618 527546 61174
rect 528102 60618 528134 61174
rect 527514 25174 528134 60618
rect 527514 24618 527546 25174
rect 528102 24618 528134 25174
rect 527514 -3226 528134 24618
rect 527514 -3782 527546 -3226
rect 528102 -3782 528134 -3226
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676338 531266 676894
rect 531822 676338 531854 676894
rect 531234 640894 531854 676338
rect 531234 640338 531266 640894
rect 531822 640338 531854 640894
rect 531234 604894 531854 640338
rect 531234 604338 531266 604894
rect 531822 604338 531854 604894
rect 531234 568894 531854 604338
rect 531234 568338 531266 568894
rect 531822 568338 531854 568894
rect 531234 532894 531854 568338
rect 531234 532338 531266 532894
rect 531822 532338 531854 532894
rect 531234 496894 531854 532338
rect 531234 496338 531266 496894
rect 531822 496338 531854 496894
rect 531234 460894 531854 496338
rect 531234 460338 531266 460894
rect 531822 460338 531854 460894
rect 531234 424894 531854 460338
rect 531234 424338 531266 424894
rect 531822 424338 531854 424894
rect 531234 388894 531854 424338
rect 531234 388338 531266 388894
rect 531822 388338 531854 388894
rect 531234 352894 531854 388338
rect 531234 352338 531266 352894
rect 531822 352338 531854 352894
rect 531234 316894 531854 352338
rect 531234 316338 531266 316894
rect 531822 316338 531854 316894
rect 531234 280894 531854 316338
rect 531234 280338 531266 280894
rect 531822 280338 531854 280894
rect 531234 244894 531854 280338
rect 531234 244338 531266 244894
rect 531822 244338 531854 244894
rect 531234 208894 531854 244338
rect 531234 208338 531266 208894
rect 531822 208338 531854 208894
rect 531234 172894 531854 208338
rect 531234 172338 531266 172894
rect 531822 172338 531854 172894
rect 531234 136894 531854 172338
rect 531234 136338 531266 136894
rect 531822 136338 531854 136894
rect 531234 100894 531854 136338
rect 531234 100338 531266 100894
rect 531822 100338 531854 100894
rect 531234 64894 531854 100338
rect 531234 64338 531266 64894
rect 531822 64338 531854 64894
rect 531234 28894 531854 64338
rect 531234 28338 531266 28894
rect 531822 28338 531854 28894
rect 531234 -5146 531854 28338
rect 531234 -5702 531266 -5146
rect 531822 -5702 531854 -5146
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710042 552986 710598
rect 553542 710042 553574 710598
rect 549234 708678 549854 709670
rect 549234 708122 549266 708678
rect 549822 708122 549854 708678
rect 545514 706758 546134 707750
rect 545514 706202 545546 706758
rect 546102 706202 546134 706758
rect 534954 680058 534986 680614
rect 535542 680058 535574 680614
rect 534954 644614 535574 680058
rect 534954 644058 534986 644614
rect 535542 644058 535574 644614
rect 534954 608614 535574 644058
rect 534954 608058 534986 608614
rect 535542 608058 535574 608614
rect 534954 572614 535574 608058
rect 534954 572058 534986 572614
rect 535542 572058 535574 572614
rect 534954 536614 535574 572058
rect 534954 536058 534986 536614
rect 535542 536058 535574 536614
rect 534954 500614 535574 536058
rect 534954 500058 534986 500614
rect 535542 500058 535574 500614
rect 534954 464614 535574 500058
rect 534954 464058 534986 464614
rect 535542 464058 535574 464614
rect 534954 428614 535574 464058
rect 534954 428058 534986 428614
rect 535542 428058 535574 428614
rect 534954 392614 535574 428058
rect 534954 392058 534986 392614
rect 535542 392058 535574 392614
rect 534954 356614 535574 392058
rect 534954 356058 534986 356614
rect 535542 356058 535574 356614
rect 534954 320614 535574 356058
rect 534954 320058 534986 320614
rect 535542 320058 535574 320614
rect 534954 284614 535574 320058
rect 534954 284058 534986 284614
rect 535542 284058 535574 284614
rect 534954 248614 535574 284058
rect 534954 248058 534986 248614
rect 535542 248058 535574 248614
rect 534954 212614 535574 248058
rect 534954 212058 534986 212614
rect 535542 212058 535574 212614
rect 534954 176614 535574 212058
rect 534954 176058 534986 176614
rect 535542 176058 535574 176614
rect 534954 140614 535574 176058
rect 534954 140058 534986 140614
rect 535542 140058 535574 140614
rect 534954 104614 535574 140058
rect 534954 104058 534986 104614
rect 535542 104058 535574 104614
rect 534954 68614 535574 104058
rect 534954 68058 534986 68614
rect 535542 68058 535574 68614
rect 534954 32614 535574 68058
rect 534954 32058 534986 32614
rect 535542 32058 535574 32614
rect 516954 -6662 516986 -6106
rect 517542 -6662 517574 -6106
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704282 541826 704838
rect 542382 704282 542414 704838
rect 541794 687454 542414 704282
rect 541794 686898 541826 687454
rect 542382 686898 542414 687454
rect 541794 651454 542414 686898
rect 541794 650898 541826 651454
rect 542382 650898 542414 651454
rect 541794 615454 542414 650898
rect 541794 614898 541826 615454
rect 542382 614898 542414 615454
rect 541794 579454 542414 614898
rect 541794 578898 541826 579454
rect 542382 578898 542414 579454
rect 541794 543454 542414 578898
rect 541794 542898 541826 543454
rect 542382 542898 542414 543454
rect 541794 507454 542414 542898
rect 541794 506898 541826 507454
rect 542382 506898 542414 507454
rect 541794 471454 542414 506898
rect 541794 470898 541826 471454
rect 542382 470898 542414 471454
rect 541794 435454 542414 470898
rect 541794 434898 541826 435454
rect 542382 434898 542414 435454
rect 541794 399454 542414 434898
rect 541794 398898 541826 399454
rect 542382 398898 542414 399454
rect 541794 363454 542414 398898
rect 541794 362898 541826 363454
rect 542382 362898 542414 363454
rect 541794 327454 542414 362898
rect 541794 326898 541826 327454
rect 542382 326898 542414 327454
rect 541794 291454 542414 326898
rect 541794 290898 541826 291454
rect 542382 290898 542414 291454
rect 541794 255454 542414 290898
rect 541794 254898 541826 255454
rect 542382 254898 542414 255454
rect 541794 219454 542414 254898
rect 541794 218898 541826 219454
rect 542382 218898 542414 219454
rect 541794 183454 542414 218898
rect 541794 182898 541826 183454
rect 542382 182898 542414 183454
rect 541794 147454 542414 182898
rect 541794 146898 541826 147454
rect 542382 146898 542414 147454
rect 541794 111454 542414 146898
rect 541794 110898 541826 111454
rect 542382 110898 542414 111454
rect 541794 75454 542414 110898
rect 541794 74898 541826 75454
rect 542382 74898 542414 75454
rect 541794 39454 542414 74898
rect 541794 38898 541826 39454
rect 542382 38898 542414 39454
rect 541794 3454 542414 38898
rect 541794 2898 541826 3454
rect 542382 2898 542414 3454
rect 541794 -346 542414 2898
rect 541794 -902 541826 -346
rect 542382 -902 542414 -346
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690618 545546 691174
rect 546102 690618 546134 691174
rect 545514 655174 546134 690618
rect 545514 654618 545546 655174
rect 546102 654618 546134 655174
rect 545514 619174 546134 654618
rect 545514 618618 545546 619174
rect 546102 618618 546134 619174
rect 545514 583174 546134 618618
rect 545514 582618 545546 583174
rect 546102 582618 546134 583174
rect 545514 547174 546134 582618
rect 545514 546618 545546 547174
rect 546102 546618 546134 547174
rect 545514 511174 546134 546618
rect 545514 510618 545546 511174
rect 546102 510618 546134 511174
rect 545514 475174 546134 510618
rect 545514 474618 545546 475174
rect 546102 474618 546134 475174
rect 545514 439174 546134 474618
rect 545514 438618 545546 439174
rect 546102 438618 546134 439174
rect 545514 403174 546134 438618
rect 545514 402618 545546 403174
rect 546102 402618 546134 403174
rect 545514 367174 546134 402618
rect 545514 366618 545546 367174
rect 546102 366618 546134 367174
rect 545514 331174 546134 366618
rect 545514 330618 545546 331174
rect 546102 330618 546134 331174
rect 545514 295174 546134 330618
rect 545514 294618 545546 295174
rect 546102 294618 546134 295174
rect 545514 259174 546134 294618
rect 545514 258618 545546 259174
rect 546102 258618 546134 259174
rect 545514 223174 546134 258618
rect 545514 222618 545546 223174
rect 546102 222618 546134 223174
rect 545514 187174 546134 222618
rect 545514 186618 545546 187174
rect 546102 186618 546134 187174
rect 545514 151174 546134 186618
rect 545514 150618 545546 151174
rect 546102 150618 546134 151174
rect 545514 115174 546134 150618
rect 545514 114618 545546 115174
rect 546102 114618 546134 115174
rect 545514 79174 546134 114618
rect 545514 78618 545546 79174
rect 546102 78618 546134 79174
rect 545514 43174 546134 78618
rect 545514 42618 545546 43174
rect 546102 42618 546134 43174
rect 545514 7174 546134 42618
rect 545514 6618 545546 7174
rect 546102 6618 546134 7174
rect 545514 -2266 546134 6618
rect 545514 -2822 545546 -2266
rect 546102 -2822 546134 -2266
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694338 549266 694894
rect 549822 694338 549854 694894
rect 549234 658894 549854 694338
rect 549234 658338 549266 658894
rect 549822 658338 549854 658894
rect 549234 622894 549854 658338
rect 549234 622338 549266 622894
rect 549822 622338 549854 622894
rect 549234 586894 549854 622338
rect 549234 586338 549266 586894
rect 549822 586338 549854 586894
rect 549234 550894 549854 586338
rect 549234 550338 549266 550894
rect 549822 550338 549854 550894
rect 549234 514894 549854 550338
rect 549234 514338 549266 514894
rect 549822 514338 549854 514894
rect 549234 478894 549854 514338
rect 549234 478338 549266 478894
rect 549822 478338 549854 478894
rect 549234 442894 549854 478338
rect 549234 442338 549266 442894
rect 549822 442338 549854 442894
rect 549234 406894 549854 442338
rect 549234 406338 549266 406894
rect 549822 406338 549854 406894
rect 549234 370894 549854 406338
rect 549234 370338 549266 370894
rect 549822 370338 549854 370894
rect 549234 334894 549854 370338
rect 549234 334338 549266 334894
rect 549822 334338 549854 334894
rect 549234 298894 549854 334338
rect 549234 298338 549266 298894
rect 549822 298338 549854 298894
rect 549234 262894 549854 298338
rect 549234 262338 549266 262894
rect 549822 262338 549854 262894
rect 549234 226894 549854 262338
rect 549234 226338 549266 226894
rect 549822 226338 549854 226894
rect 549234 190894 549854 226338
rect 549234 190338 549266 190894
rect 549822 190338 549854 190894
rect 549234 154894 549854 190338
rect 549234 154338 549266 154894
rect 549822 154338 549854 154894
rect 549234 118894 549854 154338
rect 549234 118338 549266 118894
rect 549822 118338 549854 118894
rect 549234 82894 549854 118338
rect 549234 82338 549266 82894
rect 549822 82338 549854 82894
rect 549234 46894 549854 82338
rect 549234 46338 549266 46894
rect 549822 46338 549854 46894
rect 549234 10894 549854 46338
rect 549234 10338 549266 10894
rect 549822 10338 549854 10894
rect 549234 -4186 549854 10338
rect 549234 -4742 549266 -4186
rect 549822 -4742 549854 -4186
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711002 570986 711558
rect 571542 711002 571574 711558
rect 567234 709638 567854 709670
rect 567234 709082 567266 709638
rect 567822 709082 567854 709638
rect 563514 707718 564134 707750
rect 563514 707162 563546 707718
rect 564102 707162 564134 707718
rect 552954 698058 552986 698614
rect 553542 698058 553574 698614
rect 552954 662614 553574 698058
rect 552954 662058 552986 662614
rect 553542 662058 553574 662614
rect 552954 626614 553574 662058
rect 552954 626058 552986 626614
rect 553542 626058 553574 626614
rect 552954 590614 553574 626058
rect 552954 590058 552986 590614
rect 553542 590058 553574 590614
rect 552954 554614 553574 590058
rect 552954 554058 552986 554614
rect 553542 554058 553574 554614
rect 552954 518614 553574 554058
rect 552954 518058 552986 518614
rect 553542 518058 553574 518614
rect 552954 482614 553574 518058
rect 552954 482058 552986 482614
rect 553542 482058 553574 482614
rect 552954 446614 553574 482058
rect 552954 446058 552986 446614
rect 553542 446058 553574 446614
rect 552954 410614 553574 446058
rect 552954 410058 552986 410614
rect 553542 410058 553574 410614
rect 552954 374614 553574 410058
rect 552954 374058 552986 374614
rect 553542 374058 553574 374614
rect 552954 338614 553574 374058
rect 552954 338058 552986 338614
rect 553542 338058 553574 338614
rect 552954 302614 553574 338058
rect 552954 302058 552986 302614
rect 553542 302058 553574 302614
rect 552954 266614 553574 302058
rect 552954 266058 552986 266614
rect 553542 266058 553574 266614
rect 552954 230614 553574 266058
rect 552954 230058 552986 230614
rect 553542 230058 553574 230614
rect 552954 194614 553574 230058
rect 552954 194058 552986 194614
rect 553542 194058 553574 194614
rect 552954 158614 553574 194058
rect 552954 158058 552986 158614
rect 553542 158058 553574 158614
rect 552954 122614 553574 158058
rect 552954 122058 552986 122614
rect 553542 122058 553574 122614
rect 552954 86614 553574 122058
rect 552954 86058 552986 86614
rect 553542 86058 553574 86614
rect 552954 50614 553574 86058
rect 552954 50058 552986 50614
rect 553542 50058 553574 50614
rect 552954 14614 553574 50058
rect 552954 14058 552986 14614
rect 553542 14058 553574 14614
rect 534954 -7622 534986 -7066
rect 535542 -7622 535574 -7066
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705242 559826 705798
rect 560382 705242 560414 705798
rect 559794 669454 560414 705242
rect 559794 668898 559826 669454
rect 560382 668898 560414 669454
rect 559794 633454 560414 668898
rect 559794 632898 559826 633454
rect 560382 632898 560414 633454
rect 559794 597454 560414 632898
rect 559794 596898 559826 597454
rect 560382 596898 560414 597454
rect 559794 561454 560414 596898
rect 559794 560898 559826 561454
rect 560382 560898 560414 561454
rect 559794 525454 560414 560898
rect 559794 524898 559826 525454
rect 560382 524898 560414 525454
rect 559794 489454 560414 524898
rect 559794 488898 559826 489454
rect 560382 488898 560414 489454
rect 559794 453454 560414 488898
rect 559794 452898 559826 453454
rect 560382 452898 560414 453454
rect 559794 417454 560414 452898
rect 559794 416898 559826 417454
rect 560382 416898 560414 417454
rect 559794 381454 560414 416898
rect 559794 380898 559826 381454
rect 560382 380898 560414 381454
rect 559794 345454 560414 380898
rect 559794 344898 559826 345454
rect 560382 344898 560414 345454
rect 559794 309454 560414 344898
rect 559794 308898 559826 309454
rect 560382 308898 560414 309454
rect 559794 273454 560414 308898
rect 559794 272898 559826 273454
rect 560382 272898 560414 273454
rect 559794 237454 560414 272898
rect 559794 236898 559826 237454
rect 560382 236898 560414 237454
rect 559794 201454 560414 236898
rect 559794 200898 559826 201454
rect 560382 200898 560414 201454
rect 559794 165454 560414 200898
rect 559794 164898 559826 165454
rect 560382 164898 560414 165454
rect 559794 129454 560414 164898
rect 559794 128898 559826 129454
rect 560382 128898 560414 129454
rect 559794 93454 560414 128898
rect 559794 92898 559826 93454
rect 560382 92898 560414 93454
rect 559794 57454 560414 92898
rect 559794 56898 559826 57454
rect 560382 56898 560414 57454
rect 559794 21454 560414 56898
rect 559794 20898 559826 21454
rect 560382 20898 560414 21454
rect 559794 -1306 560414 20898
rect 559794 -1862 559826 -1306
rect 560382 -1862 560414 -1306
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672618 563546 673174
rect 564102 672618 564134 673174
rect 563514 637174 564134 672618
rect 563514 636618 563546 637174
rect 564102 636618 564134 637174
rect 563514 601174 564134 636618
rect 563514 600618 563546 601174
rect 564102 600618 564134 601174
rect 563514 565174 564134 600618
rect 563514 564618 563546 565174
rect 564102 564618 564134 565174
rect 563514 529174 564134 564618
rect 563514 528618 563546 529174
rect 564102 528618 564134 529174
rect 563514 493174 564134 528618
rect 563514 492618 563546 493174
rect 564102 492618 564134 493174
rect 563514 457174 564134 492618
rect 563514 456618 563546 457174
rect 564102 456618 564134 457174
rect 563514 421174 564134 456618
rect 563514 420618 563546 421174
rect 564102 420618 564134 421174
rect 563514 385174 564134 420618
rect 563514 384618 563546 385174
rect 564102 384618 564134 385174
rect 563514 349174 564134 384618
rect 563514 348618 563546 349174
rect 564102 348618 564134 349174
rect 563514 313174 564134 348618
rect 563514 312618 563546 313174
rect 564102 312618 564134 313174
rect 563514 277174 564134 312618
rect 563514 276618 563546 277174
rect 564102 276618 564134 277174
rect 563514 241174 564134 276618
rect 563514 240618 563546 241174
rect 564102 240618 564134 241174
rect 563514 205174 564134 240618
rect 563514 204618 563546 205174
rect 564102 204618 564134 205174
rect 563514 169174 564134 204618
rect 563514 168618 563546 169174
rect 564102 168618 564134 169174
rect 563514 133174 564134 168618
rect 563514 132618 563546 133174
rect 564102 132618 564134 133174
rect 563514 97174 564134 132618
rect 563514 96618 563546 97174
rect 564102 96618 564134 97174
rect 563514 61174 564134 96618
rect 563514 60618 563546 61174
rect 564102 60618 564134 61174
rect 563514 25174 564134 60618
rect 563514 24618 563546 25174
rect 564102 24618 564134 25174
rect 563514 -3226 564134 24618
rect 563514 -3782 563546 -3226
rect 564102 -3782 564134 -3226
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676338 567266 676894
rect 567822 676338 567854 676894
rect 567234 640894 567854 676338
rect 567234 640338 567266 640894
rect 567822 640338 567854 640894
rect 567234 604894 567854 640338
rect 567234 604338 567266 604894
rect 567822 604338 567854 604894
rect 567234 568894 567854 604338
rect 567234 568338 567266 568894
rect 567822 568338 567854 568894
rect 567234 532894 567854 568338
rect 567234 532338 567266 532894
rect 567822 532338 567854 532894
rect 567234 496894 567854 532338
rect 567234 496338 567266 496894
rect 567822 496338 567854 496894
rect 567234 460894 567854 496338
rect 567234 460338 567266 460894
rect 567822 460338 567854 460894
rect 567234 424894 567854 460338
rect 567234 424338 567266 424894
rect 567822 424338 567854 424894
rect 567234 388894 567854 424338
rect 567234 388338 567266 388894
rect 567822 388338 567854 388894
rect 567234 352894 567854 388338
rect 567234 352338 567266 352894
rect 567822 352338 567854 352894
rect 567234 316894 567854 352338
rect 567234 316338 567266 316894
rect 567822 316338 567854 316894
rect 567234 280894 567854 316338
rect 567234 280338 567266 280894
rect 567822 280338 567854 280894
rect 567234 244894 567854 280338
rect 567234 244338 567266 244894
rect 567822 244338 567854 244894
rect 567234 208894 567854 244338
rect 567234 208338 567266 208894
rect 567822 208338 567854 208894
rect 567234 172894 567854 208338
rect 567234 172338 567266 172894
rect 567822 172338 567854 172894
rect 567234 136894 567854 172338
rect 567234 136338 567266 136894
rect 567822 136338 567854 136894
rect 567234 100894 567854 136338
rect 567234 100338 567266 100894
rect 567822 100338 567854 100894
rect 567234 64894 567854 100338
rect 567234 64338 567266 64894
rect 567822 64338 567854 64894
rect 567234 28894 567854 64338
rect 567234 28338 567266 28894
rect 567822 28338 567854 28894
rect 567234 -5146 567854 28338
rect 567234 -5702 567266 -5146
rect 567822 -5702 567854 -5146
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 581514 706202 581546 706758
rect 582102 706202 582134 706758
rect 570954 680058 570986 680614
rect 571542 680058 571574 680614
rect 570954 644614 571574 680058
rect 570954 644058 570986 644614
rect 571542 644058 571574 644614
rect 570954 608614 571574 644058
rect 570954 608058 570986 608614
rect 571542 608058 571574 608614
rect 570954 572614 571574 608058
rect 570954 572058 570986 572614
rect 571542 572058 571574 572614
rect 570954 536614 571574 572058
rect 570954 536058 570986 536614
rect 571542 536058 571574 536614
rect 570954 500614 571574 536058
rect 570954 500058 570986 500614
rect 571542 500058 571574 500614
rect 570954 464614 571574 500058
rect 577794 704838 578414 705830
rect 577794 704282 577826 704838
rect 578382 704282 578414 704838
rect 577794 687454 578414 704282
rect 577794 686898 577826 687454
rect 578382 686898 578414 687454
rect 577794 651454 578414 686898
rect 577794 650898 577826 651454
rect 578382 650898 578414 651454
rect 577794 615454 578414 650898
rect 577794 614898 577826 615454
rect 578382 614898 578414 615454
rect 577794 579454 578414 614898
rect 577794 578898 577826 579454
rect 578382 578898 578414 579454
rect 577794 543454 578414 578898
rect 577794 542898 577826 543454
rect 578382 542898 578414 543454
rect 577794 507454 578414 542898
rect 577794 506898 577826 507454
rect 578382 506898 578414 507454
rect 577451 498268 577517 498269
rect 577451 498204 577452 498268
rect 577516 498204 577517 498268
rect 577451 498203 577517 498204
rect 570954 464058 570986 464614
rect 571542 464058 571574 464614
rect 570954 428614 571574 464058
rect 570954 428058 570986 428614
rect 571542 428058 571574 428614
rect 570954 392614 571574 428058
rect 570954 392058 570986 392614
rect 571542 392058 571574 392614
rect 570954 356614 571574 392058
rect 570954 356058 570986 356614
rect 571542 356058 571574 356614
rect 570954 320614 571574 356058
rect 570954 320058 570986 320614
rect 571542 320058 571574 320614
rect 570954 284614 571574 320058
rect 570954 284058 570986 284614
rect 571542 284058 571574 284614
rect 570954 248614 571574 284058
rect 570954 248058 570986 248614
rect 571542 248058 571574 248614
rect 570954 212614 571574 248058
rect 570954 212058 570986 212614
rect 571542 212058 571574 212614
rect 570954 176614 571574 212058
rect 570954 176058 570986 176614
rect 571542 176058 571574 176614
rect 570954 140614 571574 176058
rect 570954 140058 570986 140614
rect 571542 140058 571574 140614
rect 570954 104614 571574 140058
rect 570954 104058 570986 104614
rect 571542 104058 571574 104614
rect 570954 68614 571574 104058
rect 570954 68058 570986 68614
rect 571542 68058 571574 68614
rect 570954 32614 571574 68058
rect 570954 32058 570986 32614
rect 571542 32058 571574 32614
rect 552954 -6662 552986 -6106
rect 553542 -6662 553574 -6106
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577454 19821 577514 498203
rect 577794 471454 578414 506898
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581514 690618 581546 691174
rect 582102 690618 582134 691174
rect 581514 655174 582134 690618
rect 581514 654618 581546 655174
rect 582102 654618 582134 655174
rect 581514 619174 582134 654618
rect 581514 618618 581546 619174
rect 582102 618618 582134 619174
rect 581514 583174 582134 618618
rect 581514 582618 581546 583174
rect 582102 582618 582134 583174
rect 581514 547174 582134 582618
rect 581514 546618 581546 547174
rect 582102 546618 582134 547174
rect 581514 511174 582134 546618
rect 581514 510618 581546 511174
rect 582102 510618 582134 511174
rect 580395 499900 580461 499901
rect 580395 499836 580396 499900
rect 580460 499836 580461 499900
rect 580395 499835 580461 499836
rect 580211 499764 580277 499765
rect 580211 499700 580212 499764
rect 580276 499700 580277 499764
rect 580211 499699 580277 499700
rect 577794 470898 577826 471454
rect 578382 470898 578414 471454
rect 577794 435454 578414 470898
rect 577794 434898 577826 435454
rect 578382 434898 578414 435454
rect 577794 399454 578414 434898
rect 577794 398898 577826 399454
rect 578382 398898 578414 399454
rect 577794 363454 578414 398898
rect 577794 362898 577826 363454
rect 578382 362898 578414 363454
rect 577794 327454 578414 362898
rect 577794 326898 577826 327454
rect 578382 326898 578414 327454
rect 577794 291454 578414 326898
rect 577794 290898 577826 291454
rect 578382 290898 578414 291454
rect 577794 255454 578414 290898
rect 577794 254898 577826 255454
rect 578382 254898 578414 255454
rect 577794 219454 578414 254898
rect 577794 218898 577826 219454
rect 578382 218898 578414 219454
rect 577794 183454 578414 218898
rect 577794 182898 577826 183454
rect 578382 182898 578414 183454
rect 577794 147454 578414 182898
rect 577794 146898 577826 147454
rect 578382 146898 578414 147454
rect 577794 111454 578414 146898
rect 577794 110898 577826 111454
rect 578382 110898 578414 111454
rect 577794 75454 578414 110898
rect 577794 74898 577826 75454
rect 578382 74898 578414 75454
rect 577794 39454 578414 74898
rect 580214 46341 580274 499699
rect 580398 86189 580458 499835
rect 580579 496908 580645 496909
rect 580579 496844 580580 496908
rect 580644 496844 580645 496908
rect 580579 496843 580645 496844
rect 580582 126037 580642 496843
rect 581514 475174 582134 510618
rect 581514 474618 581546 475174
rect 582102 474618 582134 475174
rect 581514 439174 582134 474618
rect 581514 438618 581546 439174
rect 582102 438618 582134 439174
rect 581514 403174 582134 438618
rect 581514 402618 581546 403174
rect 582102 402618 582134 403174
rect 581514 367174 582134 402618
rect 581514 366618 581546 367174
rect 582102 366618 582134 367174
rect 581514 331174 582134 366618
rect 581514 330618 581546 331174
rect 582102 330618 582134 331174
rect 581514 295174 582134 330618
rect 581514 294618 581546 295174
rect 582102 294618 582134 295174
rect 581514 259174 582134 294618
rect 581514 258618 581546 259174
rect 582102 258618 582134 259174
rect 581514 223174 582134 258618
rect 581514 222618 581546 223174
rect 582102 222618 582134 223174
rect 581514 187174 582134 222618
rect 581514 186618 581546 187174
rect 582102 186618 582134 187174
rect 581514 151174 582134 186618
rect 581514 150618 581546 151174
rect 582102 150618 582134 151174
rect 580579 126036 580645 126037
rect 580579 125972 580580 126036
rect 580644 125972 580645 126036
rect 580579 125971 580645 125972
rect 581514 115174 582134 150618
rect 581514 114618 581546 115174
rect 582102 114618 582134 115174
rect 580395 86188 580461 86189
rect 580395 86124 580396 86188
rect 580460 86124 580461 86188
rect 580395 86123 580461 86124
rect 581514 79174 582134 114618
rect 581514 78618 581546 79174
rect 582102 78618 582134 79174
rect 580211 46340 580277 46341
rect 580211 46276 580212 46340
rect 580276 46276 580277 46340
rect 580211 46275 580277 46276
rect 577794 38898 577826 39454
rect 578382 38898 578414 39454
rect 577451 19820 577517 19821
rect 577451 19756 577452 19820
rect 577516 19756 577517 19820
rect 577451 19755 577517 19756
rect 577794 3454 578414 38898
rect 577794 2898 577826 3454
rect 578382 2898 578414 3454
rect 577794 -346 578414 2898
rect 577794 -902 577826 -346
rect 578382 -902 578414 -346
rect 577794 -1894 578414 -902
rect 581514 43174 582134 78618
rect 581514 42618 581546 43174
rect 582102 42618 582134 43174
rect 581514 7174 582134 42618
rect 581514 6618 581546 7174
rect 582102 6618 582134 7174
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 687454 585930 704282
rect 585310 686898 585342 687454
rect 585898 686898 585930 687454
rect 585310 651454 585930 686898
rect 585310 650898 585342 651454
rect 585898 650898 585930 651454
rect 585310 615454 585930 650898
rect 585310 614898 585342 615454
rect 585898 614898 585930 615454
rect 585310 579454 585930 614898
rect 585310 578898 585342 579454
rect 585898 578898 585930 579454
rect 585310 543454 585930 578898
rect 585310 542898 585342 543454
rect 585898 542898 585930 543454
rect 585310 507454 585930 542898
rect 585310 506898 585342 507454
rect 585898 506898 585930 507454
rect 585310 471454 585930 506898
rect 585310 470898 585342 471454
rect 585898 470898 585930 471454
rect 585310 435454 585930 470898
rect 585310 434898 585342 435454
rect 585898 434898 585930 435454
rect 585310 399454 585930 434898
rect 585310 398898 585342 399454
rect 585898 398898 585930 399454
rect 585310 363454 585930 398898
rect 585310 362898 585342 363454
rect 585898 362898 585930 363454
rect 585310 327454 585930 362898
rect 585310 326898 585342 327454
rect 585898 326898 585930 327454
rect 585310 291454 585930 326898
rect 585310 290898 585342 291454
rect 585898 290898 585930 291454
rect 585310 255454 585930 290898
rect 585310 254898 585342 255454
rect 585898 254898 585930 255454
rect 585310 219454 585930 254898
rect 585310 218898 585342 219454
rect 585898 218898 585930 219454
rect 585310 183454 585930 218898
rect 585310 182898 585342 183454
rect 585898 182898 585930 183454
rect 585310 147454 585930 182898
rect 585310 146898 585342 147454
rect 585898 146898 585930 147454
rect 585310 111454 585930 146898
rect 585310 110898 585342 111454
rect 585898 110898 585930 111454
rect 585310 75454 585930 110898
rect 585310 74898 585342 75454
rect 585898 74898 585930 75454
rect 585310 39454 585930 74898
rect 585310 38898 585342 39454
rect 585898 38898 585930 39454
rect 585310 3454 585930 38898
rect 585310 2898 585342 3454
rect 585898 2898 585930 3454
rect 585310 -346 585930 2898
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 668898 586302 669454
rect 586858 668898 586890 669454
rect 586270 633454 586890 668898
rect 586270 632898 586302 633454
rect 586858 632898 586890 633454
rect 586270 597454 586890 632898
rect 586270 596898 586302 597454
rect 586858 596898 586890 597454
rect 586270 561454 586890 596898
rect 586270 560898 586302 561454
rect 586858 560898 586890 561454
rect 586270 525454 586890 560898
rect 586270 524898 586302 525454
rect 586858 524898 586890 525454
rect 586270 489454 586890 524898
rect 586270 488898 586302 489454
rect 586858 488898 586890 489454
rect 586270 453454 586890 488898
rect 586270 452898 586302 453454
rect 586858 452898 586890 453454
rect 586270 417454 586890 452898
rect 586270 416898 586302 417454
rect 586858 416898 586890 417454
rect 586270 381454 586890 416898
rect 586270 380898 586302 381454
rect 586858 380898 586890 381454
rect 586270 345454 586890 380898
rect 586270 344898 586302 345454
rect 586858 344898 586890 345454
rect 586270 309454 586890 344898
rect 586270 308898 586302 309454
rect 586858 308898 586890 309454
rect 586270 273454 586890 308898
rect 586270 272898 586302 273454
rect 586858 272898 586890 273454
rect 586270 237454 586890 272898
rect 586270 236898 586302 237454
rect 586858 236898 586890 237454
rect 586270 201454 586890 236898
rect 586270 200898 586302 201454
rect 586858 200898 586890 201454
rect 586270 165454 586890 200898
rect 586270 164898 586302 165454
rect 586858 164898 586890 165454
rect 586270 129454 586890 164898
rect 586270 128898 586302 129454
rect 586858 128898 586890 129454
rect 586270 93454 586890 128898
rect 586270 92898 586302 93454
rect 586858 92898 586890 93454
rect 586270 57454 586890 92898
rect 586270 56898 586302 57454
rect 586858 56898 586890 57454
rect 586270 21454 586890 56898
rect 586270 20898 586302 21454
rect 586858 20898 586890 21454
rect 586270 -1306 586890 20898
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690618 587262 691174
rect 587818 690618 587850 691174
rect 587230 655174 587850 690618
rect 587230 654618 587262 655174
rect 587818 654618 587850 655174
rect 587230 619174 587850 654618
rect 587230 618618 587262 619174
rect 587818 618618 587850 619174
rect 587230 583174 587850 618618
rect 587230 582618 587262 583174
rect 587818 582618 587850 583174
rect 587230 547174 587850 582618
rect 587230 546618 587262 547174
rect 587818 546618 587850 547174
rect 587230 511174 587850 546618
rect 587230 510618 587262 511174
rect 587818 510618 587850 511174
rect 587230 475174 587850 510618
rect 587230 474618 587262 475174
rect 587818 474618 587850 475174
rect 587230 439174 587850 474618
rect 587230 438618 587262 439174
rect 587818 438618 587850 439174
rect 587230 403174 587850 438618
rect 587230 402618 587262 403174
rect 587818 402618 587850 403174
rect 587230 367174 587850 402618
rect 587230 366618 587262 367174
rect 587818 366618 587850 367174
rect 587230 331174 587850 366618
rect 587230 330618 587262 331174
rect 587818 330618 587850 331174
rect 587230 295174 587850 330618
rect 587230 294618 587262 295174
rect 587818 294618 587850 295174
rect 587230 259174 587850 294618
rect 587230 258618 587262 259174
rect 587818 258618 587850 259174
rect 587230 223174 587850 258618
rect 587230 222618 587262 223174
rect 587818 222618 587850 223174
rect 587230 187174 587850 222618
rect 587230 186618 587262 187174
rect 587818 186618 587850 187174
rect 587230 151174 587850 186618
rect 587230 150618 587262 151174
rect 587818 150618 587850 151174
rect 587230 115174 587850 150618
rect 587230 114618 587262 115174
rect 587818 114618 587850 115174
rect 587230 79174 587850 114618
rect 587230 78618 587262 79174
rect 587818 78618 587850 79174
rect 587230 43174 587850 78618
rect 587230 42618 587262 43174
rect 587818 42618 587850 43174
rect 587230 7174 587850 42618
rect 587230 6618 587262 7174
rect 587818 6618 587850 7174
rect 581514 -2822 581546 -2266
rect 582102 -2822 582134 -2266
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672618 588222 673174
rect 588778 672618 588810 673174
rect 588190 637174 588810 672618
rect 588190 636618 588222 637174
rect 588778 636618 588810 637174
rect 588190 601174 588810 636618
rect 588190 600618 588222 601174
rect 588778 600618 588810 601174
rect 588190 565174 588810 600618
rect 588190 564618 588222 565174
rect 588778 564618 588810 565174
rect 588190 529174 588810 564618
rect 588190 528618 588222 529174
rect 588778 528618 588810 529174
rect 588190 493174 588810 528618
rect 588190 492618 588222 493174
rect 588778 492618 588810 493174
rect 588190 457174 588810 492618
rect 588190 456618 588222 457174
rect 588778 456618 588810 457174
rect 588190 421174 588810 456618
rect 588190 420618 588222 421174
rect 588778 420618 588810 421174
rect 588190 385174 588810 420618
rect 588190 384618 588222 385174
rect 588778 384618 588810 385174
rect 588190 349174 588810 384618
rect 588190 348618 588222 349174
rect 588778 348618 588810 349174
rect 588190 313174 588810 348618
rect 588190 312618 588222 313174
rect 588778 312618 588810 313174
rect 588190 277174 588810 312618
rect 588190 276618 588222 277174
rect 588778 276618 588810 277174
rect 588190 241174 588810 276618
rect 588190 240618 588222 241174
rect 588778 240618 588810 241174
rect 588190 205174 588810 240618
rect 588190 204618 588222 205174
rect 588778 204618 588810 205174
rect 588190 169174 588810 204618
rect 588190 168618 588222 169174
rect 588778 168618 588810 169174
rect 588190 133174 588810 168618
rect 588190 132618 588222 133174
rect 588778 132618 588810 133174
rect 588190 97174 588810 132618
rect 588190 96618 588222 97174
rect 588778 96618 588810 97174
rect 588190 61174 588810 96618
rect 588190 60618 588222 61174
rect 588778 60618 588810 61174
rect 588190 25174 588810 60618
rect 588190 24618 588222 25174
rect 588778 24618 588810 25174
rect 588190 -3226 588810 24618
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694338 589182 694894
rect 589738 694338 589770 694894
rect 589150 658894 589770 694338
rect 589150 658338 589182 658894
rect 589738 658338 589770 658894
rect 589150 622894 589770 658338
rect 589150 622338 589182 622894
rect 589738 622338 589770 622894
rect 589150 586894 589770 622338
rect 589150 586338 589182 586894
rect 589738 586338 589770 586894
rect 589150 550894 589770 586338
rect 589150 550338 589182 550894
rect 589738 550338 589770 550894
rect 589150 514894 589770 550338
rect 589150 514338 589182 514894
rect 589738 514338 589770 514894
rect 589150 478894 589770 514338
rect 589150 478338 589182 478894
rect 589738 478338 589770 478894
rect 589150 442894 589770 478338
rect 589150 442338 589182 442894
rect 589738 442338 589770 442894
rect 589150 406894 589770 442338
rect 589150 406338 589182 406894
rect 589738 406338 589770 406894
rect 589150 370894 589770 406338
rect 589150 370338 589182 370894
rect 589738 370338 589770 370894
rect 589150 334894 589770 370338
rect 589150 334338 589182 334894
rect 589738 334338 589770 334894
rect 589150 298894 589770 334338
rect 589150 298338 589182 298894
rect 589738 298338 589770 298894
rect 589150 262894 589770 298338
rect 589150 262338 589182 262894
rect 589738 262338 589770 262894
rect 589150 226894 589770 262338
rect 589150 226338 589182 226894
rect 589738 226338 589770 226894
rect 589150 190894 589770 226338
rect 589150 190338 589182 190894
rect 589738 190338 589770 190894
rect 589150 154894 589770 190338
rect 589150 154338 589182 154894
rect 589738 154338 589770 154894
rect 589150 118894 589770 154338
rect 589150 118338 589182 118894
rect 589738 118338 589770 118894
rect 589150 82894 589770 118338
rect 589150 82338 589182 82894
rect 589738 82338 589770 82894
rect 589150 46894 589770 82338
rect 589150 46338 589182 46894
rect 589738 46338 589770 46894
rect 589150 10894 589770 46338
rect 589150 10338 589182 10894
rect 589738 10338 589770 10894
rect 589150 -4186 589770 10338
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676338 590142 676894
rect 590698 676338 590730 676894
rect 590110 640894 590730 676338
rect 590110 640338 590142 640894
rect 590698 640338 590730 640894
rect 590110 604894 590730 640338
rect 590110 604338 590142 604894
rect 590698 604338 590730 604894
rect 590110 568894 590730 604338
rect 590110 568338 590142 568894
rect 590698 568338 590730 568894
rect 590110 532894 590730 568338
rect 590110 532338 590142 532894
rect 590698 532338 590730 532894
rect 590110 496894 590730 532338
rect 590110 496338 590142 496894
rect 590698 496338 590730 496894
rect 590110 460894 590730 496338
rect 590110 460338 590142 460894
rect 590698 460338 590730 460894
rect 590110 424894 590730 460338
rect 590110 424338 590142 424894
rect 590698 424338 590730 424894
rect 590110 388894 590730 424338
rect 590110 388338 590142 388894
rect 590698 388338 590730 388894
rect 590110 352894 590730 388338
rect 590110 352338 590142 352894
rect 590698 352338 590730 352894
rect 590110 316894 590730 352338
rect 590110 316338 590142 316894
rect 590698 316338 590730 316894
rect 590110 280894 590730 316338
rect 590110 280338 590142 280894
rect 590698 280338 590730 280894
rect 590110 244894 590730 280338
rect 590110 244338 590142 244894
rect 590698 244338 590730 244894
rect 590110 208894 590730 244338
rect 590110 208338 590142 208894
rect 590698 208338 590730 208894
rect 590110 172894 590730 208338
rect 590110 172338 590142 172894
rect 590698 172338 590730 172894
rect 590110 136894 590730 172338
rect 590110 136338 590142 136894
rect 590698 136338 590730 136894
rect 590110 100894 590730 136338
rect 590110 100338 590142 100894
rect 590698 100338 590730 100894
rect 590110 64894 590730 100338
rect 590110 64338 590142 64894
rect 590698 64338 590730 64894
rect 590110 28894 590730 64338
rect 590110 28338 590142 28894
rect 590698 28338 590730 28894
rect 590110 -5146 590730 28338
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698058 591102 698614
rect 591658 698058 591690 698614
rect 591070 662614 591690 698058
rect 591070 662058 591102 662614
rect 591658 662058 591690 662614
rect 591070 626614 591690 662058
rect 591070 626058 591102 626614
rect 591658 626058 591690 626614
rect 591070 590614 591690 626058
rect 591070 590058 591102 590614
rect 591658 590058 591690 590614
rect 591070 554614 591690 590058
rect 591070 554058 591102 554614
rect 591658 554058 591690 554614
rect 591070 518614 591690 554058
rect 591070 518058 591102 518614
rect 591658 518058 591690 518614
rect 591070 482614 591690 518058
rect 591070 482058 591102 482614
rect 591658 482058 591690 482614
rect 591070 446614 591690 482058
rect 591070 446058 591102 446614
rect 591658 446058 591690 446614
rect 591070 410614 591690 446058
rect 591070 410058 591102 410614
rect 591658 410058 591690 410614
rect 591070 374614 591690 410058
rect 591070 374058 591102 374614
rect 591658 374058 591690 374614
rect 591070 338614 591690 374058
rect 591070 338058 591102 338614
rect 591658 338058 591690 338614
rect 591070 302614 591690 338058
rect 591070 302058 591102 302614
rect 591658 302058 591690 302614
rect 591070 266614 591690 302058
rect 591070 266058 591102 266614
rect 591658 266058 591690 266614
rect 591070 230614 591690 266058
rect 591070 230058 591102 230614
rect 591658 230058 591690 230614
rect 591070 194614 591690 230058
rect 591070 194058 591102 194614
rect 591658 194058 591690 194614
rect 591070 158614 591690 194058
rect 591070 158058 591102 158614
rect 591658 158058 591690 158614
rect 591070 122614 591690 158058
rect 591070 122058 591102 122614
rect 591658 122058 591690 122614
rect 591070 86614 591690 122058
rect 591070 86058 591102 86614
rect 591658 86058 591690 86614
rect 591070 50614 591690 86058
rect 591070 50058 591102 50614
rect 591658 50058 591690 50614
rect 591070 14614 591690 50058
rect 591070 14058 591102 14614
rect 591658 14058 591690 14614
rect 591070 -6106 591690 14058
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680058 592062 680614
rect 592618 680058 592650 680614
rect 592030 644614 592650 680058
rect 592030 644058 592062 644614
rect 592618 644058 592650 644614
rect 592030 608614 592650 644058
rect 592030 608058 592062 608614
rect 592618 608058 592650 608614
rect 592030 572614 592650 608058
rect 592030 572058 592062 572614
rect 592618 572058 592650 572614
rect 592030 536614 592650 572058
rect 592030 536058 592062 536614
rect 592618 536058 592650 536614
rect 592030 500614 592650 536058
rect 592030 500058 592062 500614
rect 592618 500058 592650 500614
rect 592030 464614 592650 500058
rect 592030 464058 592062 464614
rect 592618 464058 592650 464614
rect 592030 428614 592650 464058
rect 592030 428058 592062 428614
rect 592618 428058 592650 428614
rect 592030 392614 592650 428058
rect 592030 392058 592062 392614
rect 592618 392058 592650 392614
rect 592030 356614 592650 392058
rect 592030 356058 592062 356614
rect 592618 356058 592650 356614
rect 592030 320614 592650 356058
rect 592030 320058 592062 320614
rect 592618 320058 592650 320614
rect 592030 284614 592650 320058
rect 592030 284058 592062 284614
rect 592618 284058 592650 284614
rect 592030 248614 592650 284058
rect 592030 248058 592062 248614
rect 592618 248058 592650 248614
rect 592030 212614 592650 248058
rect 592030 212058 592062 212614
rect 592618 212058 592650 212614
rect 592030 176614 592650 212058
rect 592030 176058 592062 176614
rect 592618 176058 592650 176614
rect 592030 140614 592650 176058
rect 592030 140058 592062 140614
rect 592618 140058 592650 140614
rect 592030 104614 592650 140058
rect 592030 104058 592062 104614
rect 592618 104058 592650 104614
rect 592030 68614 592650 104058
rect 592030 68058 592062 68614
rect 592618 68058 592650 68614
rect 592030 32614 592650 68058
rect 592030 32058 592062 32614
rect 592618 32058 592650 32614
rect 570954 -7622 570986 -7066
rect 571542 -7622 571574 -7066
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 680058 -8138 680614
rect -8694 644058 -8138 644614
rect -8694 608058 -8138 608614
rect -8694 572058 -8138 572614
rect -8694 536058 -8138 536614
rect -8694 500058 -8138 500614
rect -8694 464058 -8138 464614
rect -8694 428058 -8138 428614
rect -8694 392058 -8138 392614
rect -8694 356058 -8138 356614
rect -8694 320058 -8138 320614
rect -8694 284058 -8138 284614
rect -8694 248058 -8138 248614
rect -8694 212058 -8138 212614
rect -8694 176058 -8138 176614
rect -8694 140058 -8138 140614
rect -8694 104058 -8138 104614
rect -8694 68058 -8138 68614
rect -8694 32058 -8138 32614
rect -7734 710042 -7178 710598
rect 12986 710042 13542 710598
rect -7734 698058 -7178 698614
rect -7734 662058 -7178 662614
rect -7734 626058 -7178 626614
rect -7734 590058 -7178 590614
rect -7734 554058 -7178 554614
rect -7734 518058 -7178 518614
rect -7734 482058 -7178 482614
rect -7734 446058 -7178 446614
rect -7734 410058 -7178 410614
rect -7734 374058 -7178 374614
rect -7734 338058 -7178 338614
rect -7734 302058 -7178 302614
rect -7734 266058 -7178 266614
rect -7734 230058 -7178 230614
rect -7734 194058 -7178 194614
rect -7734 158058 -7178 158614
rect -7734 122058 -7178 122614
rect -7734 86058 -7178 86614
rect -7734 50058 -7178 50614
rect -7734 14058 -7178 14614
rect -6774 709082 -6218 709638
rect -6774 676338 -6218 676894
rect -6774 640338 -6218 640894
rect -6774 604338 -6218 604894
rect -6774 568338 -6218 568894
rect -6774 532338 -6218 532894
rect -6774 496338 -6218 496894
rect -6774 460338 -6218 460894
rect -6774 424338 -6218 424894
rect -6774 388338 -6218 388894
rect -6774 352338 -6218 352894
rect -6774 316338 -6218 316894
rect -6774 280338 -6218 280894
rect -6774 244338 -6218 244894
rect -6774 208338 -6218 208894
rect -6774 172338 -6218 172894
rect -6774 136338 -6218 136894
rect -6774 100338 -6218 100894
rect -6774 64338 -6218 64894
rect -6774 28338 -6218 28894
rect -5814 708122 -5258 708678
rect 9266 708122 9822 708678
rect -5814 694338 -5258 694894
rect -5814 658338 -5258 658894
rect -5814 622338 -5258 622894
rect -5814 586338 -5258 586894
rect -5814 550338 -5258 550894
rect -5814 514338 -5258 514894
rect -5814 478338 -5258 478894
rect -5814 442338 -5258 442894
rect -5814 406338 -5258 406894
rect -5814 370338 -5258 370894
rect -5814 334338 -5258 334894
rect -5814 298338 -5258 298894
rect -5814 262338 -5258 262894
rect -5814 226338 -5258 226894
rect -5814 190338 -5258 190894
rect -5814 154338 -5258 154894
rect -5814 118338 -5258 118894
rect -5814 82338 -5258 82894
rect -5814 46338 -5258 46894
rect -5814 10338 -5258 10894
rect -4854 707162 -4298 707718
rect -4854 672618 -4298 673174
rect -4854 636618 -4298 637174
rect -4854 600618 -4298 601174
rect -4854 564618 -4298 565174
rect -4854 528618 -4298 529174
rect -4854 492618 -4298 493174
rect -4854 456618 -4298 457174
rect -4854 420618 -4298 421174
rect -4854 384618 -4298 385174
rect -4854 348618 -4298 349174
rect -4854 312618 -4298 313174
rect -4854 276618 -4298 277174
rect -4854 240618 -4298 241174
rect -4854 204618 -4298 205174
rect -4854 168618 -4298 169174
rect -4854 132618 -4298 133174
rect -4854 96618 -4298 97174
rect -4854 60618 -4298 61174
rect -4854 24618 -4298 25174
rect -3894 706202 -3338 706758
rect 5546 706202 6102 706758
rect -3894 690618 -3338 691174
rect -3894 654618 -3338 655174
rect -3894 618618 -3338 619174
rect -3894 582618 -3338 583174
rect -3894 546618 -3338 547174
rect -3894 510618 -3338 511174
rect -3894 474618 -3338 475174
rect -3894 438618 -3338 439174
rect -3894 402618 -3338 403174
rect -3894 366618 -3338 367174
rect -3894 330618 -3338 331174
rect -3894 294618 -3338 295174
rect -3894 258618 -3338 259174
rect -3894 222618 -3338 223174
rect -3894 186618 -3338 187174
rect -3894 150618 -3338 151174
rect -3894 114618 -3338 115174
rect -3894 78618 -3338 79174
rect -3894 42618 -3338 43174
rect -3894 6618 -3338 7174
rect -2934 705242 -2378 705798
rect -2934 668898 -2378 669454
rect -2934 632898 -2378 633454
rect -2934 596898 -2378 597454
rect -2934 560898 -2378 561454
rect -2934 524898 -2378 525454
rect -2934 488898 -2378 489454
rect -2934 452898 -2378 453454
rect -2934 416898 -2378 417454
rect -2934 380898 -2378 381454
rect -2934 344898 -2378 345454
rect -2934 308898 -2378 309454
rect -2934 272898 -2378 273454
rect -2934 236898 -2378 237454
rect -2934 200898 -2378 201454
rect -2934 164898 -2378 165454
rect -2934 128898 -2378 129454
rect -2934 92898 -2378 93454
rect -2934 56898 -2378 57454
rect -2934 20898 -2378 21454
rect -1974 704282 -1418 704838
rect -1974 686898 -1418 687454
rect -1974 650898 -1418 651454
rect -1974 614898 -1418 615454
rect -1974 578898 -1418 579454
rect -1974 542898 -1418 543454
rect -1974 506898 -1418 507454
rect -1974 470898 -1418 471454
rect -1974 434898 -1418 435454
rect -1974 398898 -1418 399454
rect -1974 362898 -1418 363454
rect -1974 326898 -1418 327454
rect -1974 290898 -1418 291454
rect -1974 254898 -1418 255454
rect -1974 218898 -1418 219454
rect -1974 182898 -1418 183454
rect -1974 146898 -1418 147454
rect -1974 110898 -1418 111454
rect -1974 74898 -1418 75454
rect -1974 38898 -1418 39454
rect -1974 2898 -1418 3454
rect -1974 -902 -1418 -346
rect 1826 704282 2382 704838
rect 1826 686898 2382 687454
rect 1826 650898 2382 651454
rect 1826 614898 2382 615454
rect 1826 578898 2382 579454
rect 1826 542898 2382 543454
rect 1826 506898 2382 507454
rect 1826 470898 2382 471454
rect 1826 434898 2382 435454
rect 1826 398898 2382 399454
rect 1826 362898 2382 363454
rect 1826 326898 2382 327454
rect 1826 290898 2382 291454
rect 1826 254898 2382 255454
rect 1826 218898 2382 219454
rect 1826 182898 2382 183454
rect 1826 146898 2382 147454
rect 1826 110898 2382 111454
rect 1826 74898 2382 75454
rect 1826 38898 2382 39454
rect 1826 2898 2382 3454
rect 1826 -902 2382 -346
rect -2934 -1862 -2378 -1306
rect 5546 690618 6102 691174
rect 5546 654618 6102 655174
rect 5546 618618 6102 619174
rect 5546 582618 6102 583174
rect 5546 546618 6102 547174
rect 5546 510618 6102 511174
rect 5546 474618 6102 475174
rect 5546 438618 6102 439174
rect 5546 402618 6102 403174
rect 5546 366618 6102 367174
rect 5546 330618 6102 331174
rect 5546 294618 6102 295174
rect 5546 258618 6102 259174
rect 5546 222618 6102 223174
rect 5546 186618 6102 187174
rect 5546 150618 6102 151174
rect 5546 114618 6102 115174
rect 5546 78618 6102 79174
rect 5546 42618 6102 43174
rect 5546 6618 6102 7174
rect -3894 -2822 -3338 -2266
rect 5546 -2822 6102 -2266
rect -4854 -3782 -4298 -3226
rect 9266 694338 9822 694894
rect 9266 658338 9822 658894
rect 9266 622338 9822 622894
rect 9266 586338 9822 586894
rect 9266 550338 9822 550894
rect 9266 514338 9822 514894
rect 9266 478338 9822 478894
rect 9266 442338 9822 442894
rect 9266 406338 9822 406894
rect 9266 370338 9822 370894
rect 9266 334338 9822 334894
rect 9266 298338 9822 298894
rect 9266 262338 9822 262894
rect 9266 226338 9822 226894
rect 9266 190338 9822 190894
rect 9266 154338 9822 154894
rect 9266 118338 9822 118894
rect 9266 82338 9822 82894
rect 9266 46338 9822 46894
rect 9266 10338 9822 10894
rect -5814 -4742 -5258 -4186
rect 9266 -4742 9822 -4186
rect -6774 -5702 -6218 -5146
rect 30986 711002 31542 711558
rect 27266 709082 27822 709638
rect 23546 707162 24102 707718
rect 12986 698058 13542 698614
rect 12986 662058 13542 662614
rect 12986 626058 13542 626614
rect 12986 590058 13542 590614
rect 12986 554058 13542 554614
rect 12986 518058 13542 518614
rect 12986 482058 13542 482614
rect 12986 446058 13542 446614
rect 12986 410058 13542 410614
rect 12986 374058 13542 374614
rect 12986 338058 13542 338614
rect 12986 302058 13542 302614
rect 12986 266058 13542 266614
rect 12986 230058 13542 230614
rect 12986 194058 13542 194614
rect 12986 158058 13542 158614
rect 12986 122058 13542 122614
rect 12986 86058 13542 86614
rect 12986 50058 13542 50614
rect 12986 14058 13542 14614
rect -7734 -6662 -7178 -6106
rect 19826 705242 20382 705798
rect 19826 668898 20382 669454
rect 19826 632898 20382 633454
rect 19826 596898 20382 597454
rect 19826 560898 20382 561454
rect 19826 524898 20382 525454
rect 19826 488898 20382 489454
rect 19826 452898 20382 453454
rect 19826 416898 20382 417454
rect 19826 380898 20382 381454
rect 19826 344898 20382 345454
rect 19826 308898 20382 309454
rect 19826 272898 20382 273454
rect 19826 236898 20382 237454
rect 19826 200898 20382 201454
rect 19826 164898 20382 165454
rect 19826 128898 20382 129454
rect 19826 92898 20382 93454
rect 19826 56898 20382 57454
rect 19826 20898 20382 21454
rect 19826 -1862 20382 -1306
rect 23546 672618 24102 673174
rect 23546 636618 24102 637174
rect 23546 600618 24102 601174
rect 23546 564618 24102 565174
rect 23546 528618 24102 529174
rect 23546 492618 24102 493174
rect 23546 456618 24102 457174
rect 23546 420618 24102 421174
rect 23546 384618 24102 385174
rect 23546 348618 24102 349174
rect 23546 312618 24102 313174
rect 23546 276618 24102 277174
rect 23546 240618 24102 241174
rect 23546 204618 24102 205174
rect 23546 168618 24102 169174
rect 23546 132618 24102 133174
rect 23546 96618 24102 97174
rect 23546 60618 24102 61174
rect 23546 24618 24102 25174
rect 23546 -3782 24102 -3226
rect 27266 676338 27822 676894
rect 27266 640338 27822 640894
rect 27266 604338 27822 604894
rect 27266 568338 27822 568894
rect 27266 532338 27822 532894
rect 27266 496338 27822 496894
rect 27266 460338 27822 460894
rect 27266 424338 27822 424894
rect 27266 388338 27822 388894
rect 27266 352338 27822 352894
rect 27266 316338 27822 316894
rect 27266 280338 27822 280894
rect 27266 244338 27822 244894
rect 27266 208338 27822 208894
rect 27266 172338 27822 172894
rect 27266 136338 27822 136894
rect 27266 100338 27822 100894
rect 27266 64338 27822 64894
rect 27266 28338 27822 28894
rect 27266 -5702 27822 -5146
rect 48986 710042 49542 710598
rect 45266 708122 45822 708678
rect 41546 706202 42102 706758
rect 30986 680058 31542 680614
rect 30986 644058 31542 644614
rect 30986 608058 31542 608614
rect 30986 572058 31542 572614
rect 30986 536058 31542 536614
rect 30986 500058 31542 500614
rect 30986 464058 31542 464614
rect 30986 428058 31542 428614
rect 30986 392058 31542 392614
rect 30986 356058 31542 356614
rect 30986 320058 31542 320614
rect 30986 284058 31542 284614
rect 30986 248058 31542 248614
rect 30986 212058 31542 212614
rect 30986 176058 31542 176614
rect 30986 140058 31542 140614
rect 30986 104058 31542 104614
rect 30986 68058 31542 68614
rect 30986 32058 31542 32614
rect 12986 -6662 13542 -6106
rect -8694 -7622 -8138 -7066
rect 37826 704282 38382 704838
rect 37826 686898 38382 687454
rect 37826 650898 38382 651454
rect 37826 614898 38382 615454
rect 37826 578898 38382 579454
rect 37826 542898 38382 543454
rect 37826 506898 38382 507454
rect 37826 470898 38382 471454
rect 37826 434898 38382 435454
rect 37826 398898 38382 399454
rect 37826 362898 38382 363454
rect 37826 326898 38382 327454
rect 37826 290898 38382 291454
rect 37826 254898 38382 255454
rect 37826 218898 38382 219454
rect 37826 182898 38382 183454
rect 37826 146898 38382 147454
rect 37826 110898 38382 111454
rect 37826 74898 38382 75454
rect 37826 38898 38382 39454
rect 37826 2898 38382 3454
rect 37826 -902 38382 -346
rect 41546 690618 42102 691174
rect 41546 654618 42102 655174
rect 41546 618618 42102 619174
rect 41546 582618 42102 583174
rect 41546 546618 42102 547174
rect 41546 510618 42102 511174
rect 41546 474618 42102 475174
rect 41546 438618 42102 439174
rect 41546 402618 42102 403174
rect 41546 366618 42102 367174
rect 41546 330618 42102 331174
rect 41546 294618 42102 295174
rect 41546 258618 42102 259174
rect 41546 222618 42102 223174
rect 41546 186618 42102 187174
rect 41546 150618 42102 151174
rect 41546 114618 42102 115174
rect 41546 78618 42102 79174
rect 41546 42618 42102 43174
rect 41546 6618 42102 7174
rect 41546 -2822 42102 -2266
rect 45266 694338 45822 694894
rect 45266 658338 45822 658894
rect 45266 622338 45822 622894
rect 45266 586338 45822 586894
rect 45266 550338 45822 550894
rect 45266 514338 45822 514894
rect 45266 478338 45822 478894
rect 45266 442338 45822 442894
rect 45266 406338 45822 406894
rect 45266 370338 45822 370894
rect 45266 334338 45822 334894
rect 45266 298338 45822 298894
rect 45266 262338 45822 262894
rect 45266 226338 45822 226894
rect 45266 190338 45822 190894
rect 45266 154338 45822 154894
rect 45266 118338 45822 118894
rect 45266 82338 45822 82894
rect 45266 46338 45822 46894
rect 45266 10338 45822 10894
rect 45266 -4742 45822 -4186
rect 66986 711002 67542 711558
rect 63266 709082 63822 709638
rect 59546 707162 60102 707718
rect 48986 698058 49542 698614
rect 48986 662058 49542 662614
rect 48986 626058 49542 626614
rect 48986 590058 49542 590614
rect 48986 554058 49542 554614
rect 48986 518058 49542 518614
rect 48986 482058 49542 482614
rect 48986 446058 49542 446614
rect 48986 410058 49542 410614
rect 48986 374058 49542 374614
rect 48986 338058 49542 338614
rect 48986 302058 49542 302614
rect 48986 266058 49542 266614
rect 48986 230058 49542 230614
rect 48986 194058 49542 194614
rect 48986 158058 49542 158614
rect 48986 122058 49542 122614
rect 48986 86058 49542 86614
rect 48986 50058 49542 50614
rect 48986 14058 49542 14614
rect 30986 -7622 31542 -7066
rect 55826 705242 56382 705798
rect 55826 668898 56382 669454
rect 55826 632898 56382 633454
rect 55826 596898 56382 597454
rect 55826 560898 56382 561454
rect 55826 524898 56382 525454
rect 55826 488898 56382 489454
rect 55826 452898 56382 453454
rect 55826 416898 56382 417454
rect 55826 380898 56382 381454
rect 55826 344898 56382 345454
rect 55826 308898 56382 309454
rect 55826 272898 56382 273454
rect 55826 236898 56382 237454
rect 55826 200898 56382 201454
rect 55826 164898 56382 165454
rect 55826 128898 56382 129454
rect 55826 92898 56382 93454
rect 55826 56898 56382 57454
rect 55826 20898 56382 21454
rect 55826 -1862 56382 -1306
rect 59546 672618 60102 673174
rect 59546 636618 60102 637174
rect 59546 600618 60102 601174
rect 59546 564618 60102 565174
rect 59546 528618 60102 529174
rect 59546 492618 60102 493174
rect 59546 456618 60102 457174
rect 59546 420618 60102 421174
rect 59546 384618 60102 385174
rect 59546 348618 60102 349174
rect 59546 312618 60102 313174
rect 59546 276618 60102 277174
rect 59546 240618 60102 241174
rect 59546 204618 60102 205174
rect 59546 168618 60102 169174
rect 59546 132618 60102 133174
rect 59546 96618 60102 97174
rect 59546 60618 60102 61174
rect 59546 24618 60102 25174
rect 59546 -3782 60102 -3226
rect 63266 676338 63822 676894
rect 63266 640338 63822 640894
rect 63266 604338 63822 604894
rect 63266 568338 63822 568894
rect 63266 532338 63822 532894
rect 63266 496338 63822 496894
rect 63266 460338 63822 460894
rect 63266 424338 63822 424894
rect 63266 388338 63822 388894
rect 63266 352338 63822 352894
rect 63266 316338 63822 316894
rect 63266 280338 63822 280894
rect 63266 244338 63822 244894
rect 63266 208338 63822 208894
rect 63266 172338 63822 172894
rect 63266 136338 63822 136894
rect 63266 100338 63822 100894
rect 63266 64338 63822 64894
rect 63266 28338 63822 28894
rect 63266 -5702 63822 -5146
rect 84986 710042 85542 710598
rect 81266 708122 81822 708678
rect 77546 706202 78102 706758
rect 66986 680058 67542 680614
rect 66986 644058 67542 644614
rect 66986 608058 67542 608614
rect 66986 572058 67542 572614
rect 66986 536058 67542 536614
rect 66986 500058 67542 500614
rect 66986 464058 67542 464614
rect 66986 428058 67542 428614
rect 66986 392058 67542 392614
rect 66986 356058 67542 356614
rect 66986 320058 67542 320614
rect 66986 284058 67542 284614
rect 66986 248058 67542 248614
rect 66986 212058 67542 212614
rect 66986 176058 67542 176614
rect 66986 140058 67542 140614
rect 66986 104058 67542 104614
rect 66986 68058 67542 68614
rect 66986 32058 67542 32614
rect 48986 -6662 49542 -6106
rect 73826 704282 74382 704838
rect 73826 686898 74382 687454
rect 73826 650898 74382 651454
rect 73826 614898 74382 615454
rect 73826 578898 74382 579454
rect 73826 542898 74382 543454
rect 73826 506898 74382 507454
rect 73826 470898 74382 471454
rect 73826 434898 74382 435454
rect 73826 398898 74382 399454
rect 73826 362898 74382 363454
rect 73826 326898 74382 327454
rect 73826 290898 74382 291454
rect 73826 254898 74382 255454
rect 73826 218898 74382 219454
rect 73826 182898 74382 183454
rect 73826 146898 74382 147454
rect 73826 110898 74382 111454
rect 73826 74898 74382 75454
rect 73826 38898 74382 39454
rect 73826 2898 74382 3454
rect 73826 -902 74382 -346
rect 77546 690618 78102 691174
rect 77546 654618 78102 655174
rect 77546 618618 78102 619174
rect 77546 582618 78102 583174
rect 77546 546618 78102 547174
rect 77546 510618 78102 511174
rect 77546 474618 78102 475174
rect 77546 438618 78102 439174
rect 77546 402618 78102 403174
rect 77546 366618 78102 367174
rect 77546 330618 78102 331174
rect 77546 294618 78102 295174
rect 77546 258618 78102 259174
rect 77546 222618 78102 223174
rect 77546 186618 78102 187174
rect 77546 150618 78102 151174
rect 77546 114618 78102 115174
rect 77546 78618 78102 79174
rect 77546 42618 78102 43174
rect 77546 6618 78102 7174
rect 77546 -2822 78102 -2266
rect 81266 694338 81822 694894
rect 81266 658338 81822 658894
rect 81266 622338 81822 622894
rect 81266 586338 81822 586894
rect 81266 550338 81822 550894
rect 81266 514338 81822 514894
rect 81266 478338 81822 478894
rect 81266 442338 81822 442894
rect 81266 406338 81822 406894
rect 81266 370338 81822 370894
rect 81266 334338 81822 334894
rect 81266 298338 81822 298894
rect 81266 262338 81822 262894
rect 81266 226338 81822 226894
rect 81266 190338 81822 190894
rect 81266 154338 81822 154894
rect 81266 118338 81822 118894
rect 81266 82338 81822 82894
rect 81266 46338 81822 46894
rect 81266 10338 81822 10894
rect 81266 -4742 81822 -4186
rect 102986 711002 103542 711558
rect 99266 709082 99822 709638
rect 95546 707162 96102 707718
rect 84986 698058 85542 698614
rect 84986 662058 85542 662614
rect 84986 626058 85542 626614
rect 84986 590058 85542 590614
rect 84986 554058 85542 554614
rect 84986 518058 85542 518614
rect 84986 482058 85542 482614
rect 84986 446058 85542 446614
rect 84986 410058 85542 410614
rect 84986 374058 85542 374614
rect 84986 338058 85542 338614
rect 84986 302058 85542 302614
rect 84986 266058 85542 266614
rect 84986 230058 85542 230614
rect 84986 194058 85542 194614
rect 84986 158058 85542 158614
rect 84986 122058 85542 122614
rect 84986 86058 85542 86614
rect 84986 50058 85542 50614
rect 84986 14058 85542 14614
rect 66986 -7622 67542 -7066
rect 91826 705242 92382 705798
rect 91826 668898 92382 669454
rect 91826 632898 92382 633454
rect 91826 596898 92382 597454
rect 91826 560898 92382 561454
rect 91826 524898 92382 525454
rect 91826 488898 92382 489454
rect 91826 452898 92382 453454
rect 91826 416898 92382 417454
rect 91826 380898 92382 381454
rect 91826 344898 92382 345454
rect 91826 308898 92382 309454
rect 91826 272898 92382 273454
rect 91826 236898 92382 237454
rect 91826 200898 92382 201454
rect 91826 164898 92382 165454
rect 91826 128898 92382 129454
rect 91826 92898 92382 93454
rect 91826 56898 92382 57454
rect 91826 20898 92382 21454
rect 91826 -1862 92382 -1306
rect 95546 672618 96102 673174
rect 95546 636618 96102 637174
rect 95546 600618 96102 601174
rect 95546 564618 96102 565174
rect 95546 528618 96102 529174
rect 95546 492618 96102 493174
rect 95546 456618 96102 457174
rect 95546 420618 96102 421174
rect 95546 384618 96102 385174
rect 95546 348618 96102 349174
rect 95546 312618 96102 313174
rect 95546 276618 96102 277174
rect 95546 240618 96102 241174
rect 95546 204618 96102 205174
rect 95546 168618 96102 169174
rect 95546 132618 96102 133174
rect 95546 96618 96102 97174
rect 95546 60618 96102 61174
rect 95546 24618 96102 25174
rect 95546 -3782 96102 -3226
rect 99266 676338 99822 676894
rect 99266 640338 99822 640894
rect 99266 604338 99822 604894
rect 99266 568338 99822 568894
rect 99266 532338 99822 532894
rect 99266 496338 99822 496894
rect 99266 460338 99822 460894
rect 99266 424338 99822 424894
rect 99266 388338 99822 388894
rect 99266 352338 99822 352894
rect 99266 316338 99822 316894
rect 99266 280338 99822 280894
rect 99266 244338 99822 244894
rect 99266 208338 99822 208894
rect 99266 172338 99822 172894
rect 99266 136338 99822 136894
rect 99266 100338 99822 100894
rect 99266 64338 99822 64894
rect 99266 28338 99822 28894
rect 99266 -5702 99822 -5146
rect 120986 710042 121542 710598
rect 117266 708122 117822 708678
rect 113546 706202 114102 706758
rect 102986 680058 103542 680614
rect 102986 644058 103542 644614
rect 102986 608058 103542 608614
rect 102986 572058 103542 572614
rect 102986 536058 103542 536614
rect 102986 500058 103542 500614
rect 102986 464058 103542 464614
rect 102986 428058 103542 428614
rect 102986 392058 103542 392614
rect 102986 356058 103542 356614
rect 102986 320058 103542 320614
rect 102986 284058 103542 284614
rect 102986 248058 103542 248614
rect 102986 212058 103542 212614
rect 102986 176058 103542 176614
rect 102986 140058 103542 140614
rect 102986 104058 103542 104614
rect 102986 68058 103542 68614
rect 102986 32058 103542 32614
rect 84986 -6662 85542 -6106
rect 109826 704282 110382 704838
rect 109826 686898 110382 687454
rect 109826 650898 110382 651454
rect 109826 614898 110382 615454
rect 109826 578898 110382 579454
rect 109826 542898 110382 543454
rect 109826 506898 110382 507454
rect 109826 470898 110382 471454
rect 109826 434898 110382 435454
rect 109826 398898 110382 399454
rect 109826 362898 110382 363454
rect 109826 326898 110382 327454
rect 109826 290898 110382 291454
rect 109826 254898 110382 255454
rect 109826 218898 110382 219454
rect 109826 182898 110382 183454
rect 109826 146898 110382 147454
rect 109826 110898 110382 111454
rect 109826 74898 110382 75454
rect 109826 38898 110382 39454
rect 109826 2898 110382 3454
rect 109826 -902 110382 -346
rect 113546 690618 114102 691174
rect 113546 654618 114102 655174
rect 113546 618618 114102 619174
rect 113546 582618 114102 583174
rect 113546 546618 114102 547174
rect 113546 510618 114102 511174
rect 113546 474618 114102 475174
rect 113546 438618 114102 439174
rect 113546 402618 114102 403174
rect 113546 366618 114102 367174
rect 113546 330618 114102 331174
rect 113546 294618 114102 295174
rect 113546 258618 114102 259174
rect 113546 222618 114102 223174
rect 113546 186618 114102 187174
rect 113546 150618 114102 151174
rect 113546 114618 114102 115174
rect 113546 78618 114102 79174
rect 113546 42618 114102 43174
rect 113546 6618 114102 7174
rect 113546 -2822 114102 -2266
rect 117266 694338 117822 694894
rect 117266 658338 117822 658894
rect 117266 622338 117822 622894
rect 117266 586338 117822 586894
rect 117266 550338 117822 550894
rect 117266 514338 117822 514894
rect 117266 478338 117822 478894
rect 117266 442338 117822 442894
rect 117266 406338 117822 406894
rect 117266 370338 117822 370894
rect 117266 334338 117822 334894
rect 117266 298338 117822 298894
rect 117266 262338 117822 262894
rect 117266 226338 117822 226894
rect 117266 190338 117822 190894
rect 117266 154338 117822 154894
rect 117266 118338 117822 118894
rect 117266 82338 117822 82894
rect 117266 46338 117822 46894
rect 117266 10338 117822 10894
rect 117266 -4742 117822 -4186
rect 138986 711002 139542 711558
rect 135266 709082 135822 709638
rect 131546 707162 132102 707718
rect 120986 698058 121542 698614
rect 120986 662058 121542 662614
rect 120986 626058 121542 626614
rect 120986 590058 121542 590614
rect 120986 554058 121542 554614
rect 120986 518058 121542 518614
rect 120986 482058 121542 482614
rect 120986 446058 121542 446614
rect 120986 410058 121542 410614
rect 120986 374058 121542 374614
rect 120986 338058 121542 338614
rect 120986 302058 121542 302614
rect 120986 266058 121542 266614
rect 120986 230058 121542 230614
rect 120986 194058 121542 194614
rect 120986 158058 121542 158614
rect 120986 122058 121542 122614
rect 120986 86058 121542 86614
rect 120986 50058 121542 50614
rect 120986 14058 121542 14614
rect 102986 -7622 103542 -7066
rect 127826 705242 128382 705798
rect 127826 668898 128382 669454
rect 127826 632898 128382 633454
rect 127826 596898 128382 597454
rect 127826 560898 128382 561454
rect 127826 524898 128382 525454
rect 127826 488898 128382 489454
rect 127826 452898 128382 453454
rect 127826 416898 128382 417454
rect 127826 380898 128382 381454
rect 127826 344898 128382 345454
rect 127826 308898 128382 309454
rect 127826 272898 128382 273454
rect 127826 236898 128382 237454
rect 127826 200898 128382 201454
rect 127826 164898 128382 165454
rect 127826 128898 128382 129454
rect 127826 92898 128382 93454
rect 127826 56898 128382 57454
rect 127826 20898 128382 21454
rect 127826 -1862 128382 -1306
rect 131546 672618 132102 673174
rect 131546 636618 132102 637174
rect 131546 600618 132102 601174
rect 131546 564618 132102 565174
rect 131546 528618 132102 529174
rect 131546 492618 132102 493174
rect 131546 456618 132102 457174
rect 131546 420618 132102 421174
rect 131546 384618 132102 385174
rect 131546 348618 132102 349174
rect 131546 312618 132102 313174
rect 131546 276618 132102 277174
rect 131546 240618 132102 241174
rect 131546 204618 132102 205174
rect 131546 168618 132102 169174
rect 131546 132618 132102 133174
rect 131546 96618 132102 97174
rect 131546 60618 132102 61174
rect 131546 24618 132102 25174
rect 131546 -3782 132102 -3226
rect 135266 676338 135822 676894
rect 135266 640338 135822 640894
rect 135266 604338 135822 604894
rect 135266 568338 135822 568894
rect 135266 532338 135822 532894
rect 135266 496338 135822 496894
rect 135266 460338 135822 460894
rect 135266 424338 135822 424894
rect 135266 388338 135822 388894
rect 135266 352338 135822 352894
rect 135266 316338 135822 316894
rect 135266 280338 135822 280894
rect 135266 244338 135822 244894
rect 135266 208338 135822 208894
rect 135266 172338 135822 172894
rect 135266 136338 135822 136894
rect 135266 100338 135822 100894
rect 135266 64338 135822 64894
rect 135266 28338 135822 28894
rect 135266 -5702 135822 -5146
rect 156986 710042 157542 710598
rect 153266 708122 153822 708678
rect 149546 706202 150102 706758
rect 138986 680058 139542 680614
rect 138986 644058 139542 644614
rect 138986 608058 139542 608614
rect 138986 572058 139542 572614
rect 138986 536058 139542 536614
rect 138986 500058 139542 500614
rect 138986 464058 139542 464614
rect 138986 428058 139542 428614
rect 138986 392058 139542 392614
rect 138986 356058 139542 356614
rect 138986 320058 139542 320614
rect 138986 284058 139542 284614
rect 138986 248058 139542 248614
rect 138986 212058 139542 212614
rect 138986 176058 139542 176614
rect 138986 140058 139542 140614
rect 138986 104058 139542 104614
rect 138986 68058 139542 68614
rect 138986 32058 139542 32614
rect 120986 -6662 121542 -6106
rect 145826 704282 146382 704838
rect 145826 686898 146382 687454
rect 145826 650898 146382 651454
rect 145826 614898 146382 615454
rect 145826 578898 146382 579454
rect 145826 542898 146382 543454
rect 145826 506898 146382 507454
rect 145826 470898 146382 471454
rect 145826 434898 146382 435454
rect 145826 398898 146382 399454
rect 145826 362898 146382 363454
rect 145826 326898 146382 327454
rect 145826 290898 146382 291454
rect 145826 254898 146382 255454
rect 145826 218898 146382 219454
rect 145826 182898 146382 183454
rect 145826 146898 146382 147454
rect 145826 110898 146382 111454
rect 145826 74898 146382 75454
rect 145826 38898 146382 39454
rect 145826 2898 146382 3454
rect 145826 -902 146382 -346
rect 149546 690618 150102 691174
rect 149546 654618 150102 655174
rect 149546 618618 150102 619174
rect 149546 582618 150102 583174
rect 149546 546618 150102 547174
rect 149546 510618 150102 511174
rect 149546 474618 150102 475174
rect 149546 438618 150102 439174
rect 149546 402618 150102 403174
rect 149546 366618 150102 367174
rect 149546 330618 150102 331174
rect 149546 294618 150102 295174
rect 149546 258618 150102 259174
rect 149546 222618 150102 223174
rect 149546 186618 150102 187174
rect 149546 150618 150102 151174
rect 149546 114618 150102 115174
rect 149546 78618 150102 79174
rect 149546 42618 150102 43174
rect 149546 6618 150102 7174
rect 149546 -2822 150102 -2266
rect 153266 694338 153822 694894
rect 153266 658338 153822 658894
rect 153266 622338 153822 622894
rect 153266 586338 153822 586894
rect 153266 550338 153822 550894
rect 153266 514338 153822 514894
rect 153266 478338 153822 478894
rect 153266 442338 153822 442894
rect 153266 406338 153822 406894
rect 153266 370338 153822 370894
rect 153266 334338 153822 334894
rect 153266 298338 153822 298894
rect 153266 262338 153822 262894
rect 153266 226338 153822 226894
rect 153266 190338 153822 190894
rect 153266 154338 153822 154894
rect 153266 118338 153822 118894
rect 153266 82338 153822 82894
rect 153266 46338 153822 46894
rect 153266 10338 153822 10894
rect 153266 -4742 153822 -4186
rect 174986 711002 175542 711558
rect 171266 709082 171822 709638
rect 167546 707162 168102 707718
rect 156986 698058 157542 698614
rect 156986 662058 157542 662614
rect 156986 626058 157542 626614
rect 156986 590058 157542 590614
rect 156986 554058 157542 554614
rect 156986 518058 157542 518614
rect 156986 482058 157542 482614
rect 156986 446058 157542 446614
rect 156986 410058 157542 410614
rect 156986 374058 157542 374614
rect 156986 338058 157542 338614
rect 156986 302058 157542 302614
rect 156986 266058 157542 266614
rect 156986 230058 157542 230614
rect 156986 194058 157542 194614
rect 156986 158058 157542 158614
rect 156986 122058 157542 122614
rect 156986 86058 157542 86614
rect 156986 50058 157542 50614
rect 156986 14058 157542 14614
rect 138986 -7622 139542 -7066
rect 163826 705242 164382 705798
rect 163826 668898 164382 669454
rect 163826 632898 164382 633454
rect 163826 596898 164382 597454
rect 163826 560898 164382 561454
rect 163826 524898 164382 525454
rect 163826 488898 164382 489454
rect 163826 452898 164382 453454
rect 163826 416898 164382 417454
rect 163826 380898 164382 381454
rect 163826 344898 164382 345454
rect 163826 308898 164382 309454
rect 163826 272898 164382 273454
rect 163826 236898 164382 237454
rect 163826 200898 164382 201454
rect 163826 164898 164382 165454
rect 163826 128898 164382 129454
rect 163826 92898 164382 93454
rect 163826 56898 164382 57454
rect 163826 20898 164382 21454
rect 163826 -1862 164382 -1306
rect 167546 672618 168102 673174
rect 167546 636618 168102 637174
rect 167546 600618 168102 601174
rect 167546 564618 168102 565174
rect 167546 528618 168102 529174
rect 167546 492618 168102 493174
rect 167546 456618 168102 457174
rect 167546 420618 168102 421174
rect 167546 384618 168102 385174
rect 167546 348618 168102 349174
rect 167546 312618 168102 313174
rect 167546 276618 168102 277174
rect 167546 240618 168102 241174
rect 167546 204618 168102 205174
rect 167546 168618 168102 169174
rect 167546 132618 168102 133174
rect 167546 96618 168102 97174
rect 167546 60618 168102 61174
rect 167546 24618 168102 25174
rect 167546 -3782 168102 -3226
rect 171266 676338 171822 676894
rect 171266 640338 171822 640894
rect 171266 604338 171822 604894
rect 171266 568338 171822 568894
rect 171266 532338 171822 532894
rect 171266 496338 171822 496894
rect 171266 460338 171822 460894
rect 171266 424338 171822 424894
rect 171266 388338 171822 388894
rect 171266 352338 171822 352894
rect 171266 316338 171822 316894
rect 171266 280338 171822 280894
rect 171266 244338 171822 244894
rect 171266 208338 171822 208894
rect 171266 172338 171822 172894
rect 171266 136338 171822 136894
rect 171266 100338 171822 100894
rect 171266 64338 171822 64894
rect 171266 28338 171822 28894
rect 171266 -5702 171822 -5146
rect 192986 710042 193542 710598
rect 189266 708122 189822 708678
rect 185546 706202 186102 706758
rect 174986 680058 175542 680614
rect 174986 644058 175542 644614
rect 174986 608058 175542 608614
rect 174986 572058 175542 572614
rect 174986 536058 175542 536614
rect 174986 500058 175542 500614
rect 174986 464058 175542 464614
rect 174986 428058 175542 428614
rect 174986 392058 175542 392614
rect 174986 356058 175542 356614
rect 174986 320058 175542 320614
rect 174986 284058 175542 284614
rect 174986 248058 175542 248614
rect 174986 212058 175542 212614
rect 174986 176058 175542 176614
rect 174986 140058 175542 140614
rect 174986 104058 175542 104614
rect 174986 68058 175542 68614
rect 174986 32058 175542 32614
rect 156986 -6662 157542 -6106
rect 181826 704282 182382 704838
rect 181826 686898 182382 687454
rect 181826 650898 182382 651454
rect 181826 614898 182382 615454
rect 181826 578898 182382 579454
rect 181826 542898 182382 543454
rect 181826 506898 182382 507454
rect 181826 470898 182382 471454
rect 181826 434898 182382 435454
rect 181826 398898 182382 399454
rect 181826 362898 182382 363454
rect 181826 326898 182382 327454
rect 181826 290898 182382 291454
rect 181826 254898 182382 255454
rect 181826 218898 182382 219454
rect 181826 182898 182382 183454
rect 181826 146898 182382 147454
rect 181826 110898 182382 111454
rect 181826 74898 182382 75454
rect 181826 38898 182382 39454
rect 181826 2898 182382 3454
rect 181826 -902 182382 -346
rect 185546 690618 186102 691174
rect 185546 654618 186102 655174
rect 185546 618618 186102 619174
rect 185546 582618 186102 583174
rect 185546 546618 186102 547174
rect 185546 510618 186102 511174
rect 185546 474618 186102 475174
rect 185546 438618 186102 439174
rect 185546 402618 186102 403174
rect 185546 366618 186102 367174
rect 185546 330618 186102 331174
rect 185546 294618 186102 295174
rect 185546 258618 186102 259174
rect 185546 222618 186102 223174
rect 185546 186618 186102 187174
rect 185546 150618 186102 151174
rect 185546 114618 186102 115174
rect 185546 78618 186102 79174
rect 185546 42618 186102 43174
rect 185546 6618 186102 7174
rect 185546 -2822 186102 -2266
rect 189266 694338 189822 694894
rect 189266 658338 189822 658894
rect 189266 622338 189822 622894
rect 189266 586338 189822 586894
rect 189266 550338 189822 550894
rect 189266 514338 189822 514894
rect 189266 478338 189822 478894
rect 189266 442338 189822 442894
rect 189266 406338 189822 406894
rect 189266 370338 189822 370894
rect 189266 334338 189822 334894
rect 189266 298338 189822 298894
rect 189266 262338 189822 262894
rect 189266 226338 189822 226894
rect 189266 190338 189822 190894
rect 189266 154338 189822 154894
rect 189266 118338 189822 118894
rect 189266 82338 189822 82894
rect 189266 46338 189822 46894
rect 189266 10338 189822 10894
rect 189266 -4742 189822 -4186
rect 210986 711002 211542 711558
rect 207266 709082 207822 709638
rect 203546 707162 204102 707718
rect 192986 698058 193542 698614
rect 192986 662058 193542 662614
rect 192986 626058 193542 626614
rect 192986 590058 193542 590614
rect 192986 554058 193542 554614
rect 192986 518058 193542 518614
rect 192986 482058 193542 482614
rect 192986 446058 193542 446614
rect 192986 410058 193542 410614
rect 192986 374058 193542 374614
rect 192986 338058 193542 338614
rect 192986 302058 193542 302614
rect 192986 266058 193542 266614
rect 192986 230058 193542 230614
rect 192986 194058 193542 194614
rect 192986 158058 193542 158614
rect 192986 122058 193542 122614
rect 192986 86058 193542 86614
rect 192986 50058 193542 50614
rect 192986 14058 193542 14614
rect 174986 -7622 175542 -7066
rect 199826 705242 200382 705798
rect 199826 668898 200382 669454
rect 199826 632898 200382 633454
rect 199826 596898 200382 597454
rect 199826 560898 200382 561454
rect 199826 524898 200382 525454
rect 199826 488898 200382 489454
rect 199826 452898 200382 453454
rect 199826 416898 200382 417454
rect 199826 380898 200382 381454
rect 199826 344898 200382 345454
rect 199826 308898 200382 309454
rect 199826 272898 200382 273454
rect 199826 236898 200382 237454
rect 199826 200898 200382 201454
rect 199826 164898 200382 165454
rect 199826 128898 200382 129454
rect 199826 92898 200382 93454
rect 199826 56898 200382 57454
rect 199826 20898 200382 21454
rect 199826 -1862 200382 -1306
rect 203546 672618 204102 673174
rect 203546 636618 204102 637174
rect 203546 600618 204102 601174
rect 203546 564618 204102 565174
rect 203546 528618 204102 529174
rect 203546 492618 204102 493174
rect 203546 456618 204102 457174
rect 203546 420618 204102 421174
rect 203546 384618 204102 385174
rect 203546 348618 204102 349174
rect 203546 312618 204102 313174
rect 203546 276618 204102 277174
rect 203546 240618 204102 241174
rect 203546 204618 204102 205174
rect 203546 168618 204102 169174
rect 203546 132618 204102 133174
rect 203546 96618 204102 97174
rect 203546 60618 204102 61174
rect 203546 24618 204102 25174
rect 203546 -3782 204102 -3226
rect 207266 676338 207822 676894
rect 207266 640338 207822 640894
rect 207266 604338 207822 604894
rect 207266 568338 207822 568894
rect 207266 532338 207822 532894
rect 207266 496338 207822 496894
rect 207266 460338 207822 460894
rect 207266 424338 207822 424894
rect 207266 388338 207822 388894
rect 207266 352338 207822 352894
rect 207266 316338 207822 316894
rect 207266 280338 207822 280894
rect 207266 244338 207822 244894
rect 207266 208338 207822 208894
rect 207266 172338 207822 172894
rect 207266 136338 207822 136894
rect 207266 100338 207822 100894
rect 207266 64338 207822 64894
rect 207266 28338 207822 28894
rect 207266 -5702 207822 -5146
rect 228986 710042 229542 710598
rect 225266 708122 225822 708678
rect 221546 706202 222102 706758
rect 210986 680058 211542 680614
rect 210986 644058 211542 644614
rect 210986 608058 211542 608614
rect 210986 572058 211542 572614
rect 210986 536058 211542 536614
rect 210986 500058 211542 500614
rect 210986 464058 211542 464614
rect 210986 428058 211542 428614
rect 210986 392058 211542 392614
rect 210986 356058 211542 356614
rect 210986 320058 211542 320614
rect 210986 284058 211542 284614
rect 210986 248058 211542 248614
rect 210986 212058 211542 212614
rect 210986 176058 211542 176614
rect 210986 140058 211542 140614
rect 210986 104058 211542 104614
rect 210986 68058 211542 68614
rect 210986 32058 211542 32614
rect 192986 -6662 193542 -6106
rect 217826 704282 218382 704838
rect 217826 686898 218382 687454
rect 217826 650898 218382 651454
rect 217826 614898 218382 615454
rect 217826 578898 218382 579454
rect 217826 542898 218382 543454
rect 217826 506898 218382 507454
rect 217826 470898 218382 471454
rect 217826 434898 218382 435454
rect 217826 398898 218382 399454
rect 217826 362898 218382 363454
rect 217826 326898 218382 327454
rect 217826 290898 218382 291454
rect 217826 254898 218382 255454
rect 217826 218898 218382 219454
rect 217826 182898 218382 183454
rect 217826 146898 218382 147454
rect 217826 110898 218382 111454
rect 217826 74898 218382 75454
rect 217826 38898 218382 39454
rect 217826 2898 218382 3454
rect 217826 -902 218382 -346
rect 221546 690618 222102 691174
rect 221546 654618 222102 655174
rect 221546 618618 222102 619174
rect 221546 582618 222102 583174
rect 221546 546618 222102 547174
rect 221546 510618 222102 511174
rect 221546 474618 222102 475174
rect 221546 438618 222102 439174
rect 221546 402618 222102 403174
rect 221546 366618 222102 367174
rect 221546 330618 222102 331174
rect 221546 294618 222102 295174
rect 221546 258618 222102 259174
rect 221546 222618 222102 223174
rect 221546 186618 222102 187174
rect 221546 150618 222102 151174
rect 221546 114618 222102 115174
rect 221546 78618 222102 79174
rect 221546 42618 222102 43174
rect 221546 6618 222102 7174
rect 221546 -2822 222102 -2266
rect 225266 694338 225822 694894
rect 225266 658338 225822 658894
rect 225266 622338 225822 622894
rect 225266 586338 225822 586894
rect 225266 550338 225822 550894
rect 225266 514338 225822 514894
rect 225266 478338 225822 478894
rect 225266 442338 225822 442894
rect 225266 406338 225822 406894
rect 225266 370338 225822 370894
rect 225266 334338 225822 334894
rect 225266 298338 225822 298894
rect 225266 262338 225822 262894
rect 225266 226338 225822 226894
rect 225266 190338 225822 190894
rect 225266 154338 225822 154894
rect 225266 118338 225822 118894
rect 225266 82338 225822 82894
rect 225266 46338 225822 46894
rect 225266 10338 225822 10894
rect 225266 -4742 225822 -4186
rect 246986 711002 247542 711558
rect 243266 709082 243822 709638
rect 239546 707162 240102 707718
rect 228986 698058 229542 698614
rect 228986 662058 229542 662614
rect 228986 626058 229542 626614
rect 228986 590058 229542 590614
rect 228986 554058 229542 554614
rect 228986 518058 229542 518614
rect 235826 705242 236382 705798
rect 235826 668898 236382 669454
rect 235826 632898 236382 633454
rect 235826 596898 236382 597454
rect 235826 560898 236382 561454
rect 235826 524898 236382 525454
rect 239546 672618 240102 673174
rect 239546 636618 240102 637174
rect 239546 600618 240102 601174
rect 239546 564618 240102 565174
rect 239546 528618 240102 529174
rect 228986 482058 229542 482614
rect 228986 446058 229542 446614
rect 228986 410058 229542 410614
rect 228986 374058 229542 374614
rect 228986 338058 229542 338614
rect 228986 302058 229542 302614
rect 228986 266058 229542 266614
rect 228986 230058 229542 230614
rect 228986 194058 229542 194614
rect 228986 158058 229542 158614
rect 228986 122058 229542 122614
rect 228986 86058 229542 86614
rect 235826 308898 236382 309454
rect 235826 272898 236382 273454
rect 243266 676338 243822 676894
rect 243266 640338 243822 640894
rect 243266 604338 243822 604894
rect 243266 568338 243822 568894
rect 243266 532338 243822 532894
rect 264986 710042 265542 710598
rect 261266 708122 261822 708678
rect 257546 706202 258102 706758
rect 246986 680058 247542 680614
rect 246986 644058 247542 644614
rect 246986 608058 247542 608614
rect 246986 572058 247542 572614
rect 246986 536058 247542 536614
rect 246986 500058 247542 500614
rect 253826 704282 254382 704838
rect 253826 686898 254382 687454
rect 253826 650898 254382 651454
rect 253826 614898 254382 615454
rect 253826 578898 254382 579454
rect 253826 542898 254382 543454
rect 253826 506898 254382 507454
rect 257546 690618 258102 691174
rect 257546 654618 258102 655174
rect 257546 618618 258102 619174
rect 257546 582618 258102 583174
rect 257546 546618 258102 547174
rect 257546 510618 258102 511174
rect 261266 694338 261822 694894
rect 261266 658338 261822 658894
rect 261266 622338 261822 622894
rect 261266 586338 261822 586894
rect 261266 550338 261822 550894
rect 261266 514338 261822 514894
rect 282986 711002 283542 711558
rect 279266 709082 279822 709638
rect 275546 707162 276102 707718
rect 264986 698058 265542 698614
rect 264986 662058 265542 662614
rect 264986 626058 265542 626614
rect 264986 590058 265542 590614
rect 264986 554058 265542 554614
rect 264986 518058 265542 518614
rect 271826 705242 272382 705798
rect 271826 668898 272382 669454
rect 271826 632898 272382 633454
rect 271826 596898 272382 597454
rect 271826 560898 272382 561454
rect 271826 524898 272382 525454
rect 275546 672618 276102 673174
rect 275546 636618 276102 637174
rect 275546 600618 276102 601174
rect 275546 564618 276102 565174
rect 275546 528618 276102 529174
rect 279266 676338 279822 676894
rect 279266 640338 279822 640894
rect 279266 604338 279822 604894
rect 279266 568338 279822 568894
rect 279266 532338 279822 532894
rect 300986 710042 301542 710598
rect 297266 708122 297822 708678
rect 293546 706202 294102 706758
rect 282986 680058 283542 680614
rect 282986 644058 283542 644614
rect 282986 608058 283542 608614
rect 282986 572058 283542 572614
rect 282986 536058 283542 536614
rect 282986 500058 283542 500614
rect 289826 704282 290382 704838
rect 289826 686898 290382 687454
rect 289826 650898 290382 651454
rect 289826 614898 290382 615454
rect 289826 578898 290382 579454
rect 289826 542898 290382 543454
rect 289826 506898 290382 507454
rect 293546 690618 294102 691174
rect 293546 654618 294102 655174
rect 293546 618618 294102 619174
rect 293546 582618 294102 583174
rect 293546 546618 294102 547174
rect 293546 510618 294102 511174
rect 297266 694338 297822 694894
rect 297266 658338 297822 658894
rect 297266 622338 297822 622894
rect 297266 586338 297822 586894
rect 297266 550338 297822 550894
rect 297266 514338 297822 514894
rect 318986 711002 319542 711558
rect 315266 709082 315822 709638
rect 311546 707162 312102 707718
rect 300986 698058 301542 698614
rect 300986 662058 301542 662614
rect 300986 626058 301542 626614
rect 300986 590058 301542 590614
rect 300986 554058 301542 554614
rect 300986 518058 301542 518614
rect 307826 705242 308382 705798
rect 307826 668898 308382 669454
rect 307826 632898 308382 633454
rect 307826 596898 308382 597454
rect 307826 560898 308382 561454
rect 307826 524898 308382 525454
rect 311546 672618 312102 673174
rect 311546 636618 312102 637174
rect 311546 600618 312102 601174
rect 311546 564618 312102 565174
rect 311546 528618 312102 529174
rect 315266 676338 315822 676894
rect 315266 640338 315822 640894
rect 315266 604338 315822 604894
rect 315266 568338 315822 568894
rect 315266 532338 315822 532894
rect 336986 710042 337542 710598
rect 333266 708122 333822 708678
rect 329546 706202 330102 706758
rect 318986 680058 319542 680614
rect 318986 644058 319542 644614
rect 318986 608058 319542 608614
rect 318986 572058 319542 572614
rect 318986 536058 319542 536614
rect 318986 500058 319542 500614
rect 325826 704282 326382 704838
rect 325826 686898 326382 687454
rect 325826 650898 326382 651454
rect 325826 614898 326382 615454
rect 325826 578898 326382 579454
rect 325826 542898 326382 543454
rect 325826 506898 326382 507454
rect 329546 690618 330102 691174
rect 329546 654618 330102 655174
rect 329546 618618 330102 619174
rect 329546 582618 330102 583174
rect 329546 546618 330102 547174
rect 329546 510618 330102 511174
rect 333266 694338 333822 694894
rect 333266 658338 333822 658894
rect 333266 622338 333822 622894
rect 333266 586338 333822 586894
rect 333266 550338 333822 550894
rect 333266 514338 333822 514894
rect 354986 711002 355542 711558
rect 351266 709082 351822 709638
rect 347546 707162 348102 707718
rect 336986 698058 337542 698614
rect 336986 662058 337542 662614
rect 336986 626058 337542 626614
rect 336986 590058 337542 590614
rect 336986 554058 337542 554614
rect 336986 518058 337542 518614
rect 343826 705242 344382 705798
rect 343826 668898 344382 669454
rect 343826 632898 344382 633454
rect 343826 596898 344382 597454
rect 343826 560898 344382 561454
rect 343826 524898 344382 525454
rect 347546 672618 348102 673174
rect 347546 636618 348102 637174
rect 347546 600618 348102 601174
rect 347546 564618 348102 565174
rect 347546 528618 348102 529174
rect 351266 676338 351822 676894
rect 351266 640338 351822 640894
rect 351266 604338 351822 604894
rect 351266 568338 351822 568894
rect 351266 532338 351822 532894
rect 372986 710042 373542 710598
rect 369266 708122 369822 708678
rect 365546 706202 366102 706758
rect 354986 680058 355542 680614
rect 354986 644058 355542 644614
rect 354986 608058 355542 608614
rect 354986 572058 355542 572614
rect 354986 536058 355542 536614
rect 354986 500058 355542 500614
rect 361826 704282 362382 704838
rect 361826 686898 362382 687454
rect 361826 650898 362382 651454
rect 361826 614898 362382 615454
rect 361826 578898 362382 579454
rect 361826 542898 362382 543454
rect 361826 506898 362382 507454
rect 365546 690618 366102 691174
rect 365546 654618 366102 655174
rect 365546 618618 366102 619174
rect 365546 582618 366102 583174
rect 365546 546618 366102 547174
rect 365546 510618 366102 511174
rect 369266 694338 369822 694894
rect 369266 658338 369822 658894
rect 369266 622338 369822 622894
rect 369266 586338 369822 586894
rect 369266 550338 369822 550894
rect 369266 514338 369822 514894
rect 390986 711002 391542 711558
rect 387266 709082 387822 709638
rect 383546 707162 384102 707718
rect 372986 698058 373542 698614
rect 372986 662058 373542 662614
rect 372986 626058 373542 626614
rect 372986 590058 373542 590614
rect 372986 554058 373542 554614
rect 372986 518058 373542 518614
rect 379826 705242 380382 705798
rect 379826 668898 380382 669454
rect 379826 632898 380382 633454
rect 379826 596898 380382 597454
rect 379826 560898 380382 561454
rect 379826 524898 380382 525454
rect 383546 672618 384102 673174
rect 383546 636618 384102 637174
rect 383546 600618 384102 601174
rect 383546 564618 384102 565174
rect 383546 528618 384102 529174
rect 387266 676338 387822 676894
rect 387266 640338 387822 640894
rect 387266 604338 387822 604894
rect 387266 568338 387822 568894
rect 387266 532338 387822 532894
rect 408986 710042 409542 710598
rect 405266 708122 405822 708678
rect 401546 706202 402102 706758
rect 390986 680058 391542 680614
rect 390986 644058 391542 644614
rect 390986 608058 391542 608614
rect 390986 572058 391542 572614
rect 390986 536058 391542 536614
rect 390986 500058 391542 500614
rect 397826 704282 398382 704838
rect 397826 686898 398382 687454
rect 397826 650898 398382 651454
rect 397826 614898 398382 615454
rect 397826 578898 398382 579454
rect 397826 542898 398382 543454
rect 397826 506898 398382 507454
rect 401546 690618 402102 691174
rect 401546 654618 402102 655174
rect 401546 618618 402102 619174
rect 401546 582618 402102 583174
rect 401546 546618 402102 547174
rect 401546 510618 402102 511174
rect 405266 694338 405822 694894
rect 405266 658338 405822 658894
rect 405266 622338 405822 622894
rect 405266 586338 405822 586894
rect 405266 550338 405822 550894
rect 405266 514338 405822 514894
rect 426986 711002 427542 711558
rect 423266 709082 423822 709638
rect 419546 707162 420102 707718
rect 408986 698058 409542 698614
rect 408986 662058 409542 662614
rect 408986 626058 409542 626614
rect 408986 590058 409542 590614
rect 408986 554058 409542 554614
rect 408986 518058 409542 518614
rect 415826 705242 416382 705798
rect 415826 668898 416382 669454
rect 415826 632898 416382 633454
rect 415826 596898 416382 597454
rect 415826 560898 416382 561454
rect 415826 524898 416382 525454
rect 419546 672618 420102 673174
rect 419546 636618 420102 637174
rect 419546 600618 420102 601174
rect 419546 564618 420102 565174
rect 419546 528618 420102 529174
rect 423266 676338 423822 676894
rect 423266 640338 423822 640894
rect 423266 604338 423822 604894
rect 423266 568338 423822 568894
rect 423266 532338 423822 532894
rect 444986 710042 445542 710598
rect 441266 708122 441822 708678
rect 437546 706202 438102 706758
rect 426986 680058 427542 680614
rect 426986 644058 427542 644614
rect 426986 608058 427542 608614
rect 426986 572058 427542 572614
rect 426986 536058 427542 536614
rect 426986 500058 427542 500614
rect 433826 704282 434382 704838
rect 433826 686898 434382 687454
rect 433826 650898 434382 651454
rect 433826 614898 434382 615454
rect 433826 578898 434382 579454
rect 433826 542898 434382 543454
rect 433826 506898 434382 507454
rect 437546 690618 438102 691174
rect 437546 654618 438102 655174
rect 437546 618618 438102 619174
rect 437546 582618 438102 583174
rect 437546 546618 438102 547174
rect 437546 510618 438102 511174
rect 235826 236898 236382 237454
rect 235826 200898 236382 201454
rect 235826 164898 236382 165454
rect 235826 128898 236382 129454
rect 235826 92898 236382 93454
rect 228986 50058 229542 50614
rect 228986 14058 229542 14614
rect 210986 -7622 211542 -7066
rect 235826 56898 236382 57454
rect 254610 489218 254846 489454
rect 254610 488898 254846 489134
rect 285330 489218 285566 489454
rect 285330 488898 285566 489134
rect 316050 489218 316286 489454
rect 316050 488898 316286 489134
rect 346770 489218 347006 489454
rect 346770 488898 347006 489134
rect 377490 489218 377726 489454
rect 377490 488898 377726 489134
rect 408210 489218 408446 489454
rect 408210 488898 408446 489134
rect 239250 471218 239486 471454
rect 239250 470898 239486 471134
rect 269970 471218 270206 471454
rect 269970 470898 270206 471134
rect 300690 471218 300926 471454
rect 300690 470898 300926 471134
rect 331410 471218 331646 471454
rect 331410 470898 331646 471134
rect 362130 471218 362366 471454
rect 362130 470898 362366 471134
rect 392850 471218 393086 471454
rect 392850 470898 393086 471134
rect 423570 471218 423806 471454
rect 423570 470898 423806 471134
rect 254610 453218 254846 453454
rect 254610 452898 254846 453134
rect 285330 453218 285566 453454
rect 285330 452898 285566 453134
rect 316050 453218 316286 453454
rect 316050 452898 316286 453134
rect 346770 453218 347006 453454
rect 346770 452898 347006 453134
rect 377490 453218 377726 453454
rect 377490 452898 377726 453134
rect 408210 453218 408446 453454
rect 408210 452898 408446 453134
rect 239250 435218 239486 435454
rect 239250 434898 239486 435134
rect 269970 435218 270206 435454
rect 269970 434898 270206 435134
rect 300690 435218 300926 435454
rect 300690 434898 300926 435134
rect 331410 435218 331646 435454
rect 331410 434898 331646 435134
rect 362130 435218 362366 435454
rect 362130 434898 362366 435134
rect 392850 435218 393086 435454
rect 392850 434898 393086 435134
rect 423570 435218 423806 435454
rect 423570 434898 423806 435134
rect 254610 417218 254846 417454
rect 254610 416898 254846 417134
rect 285330 417218 285566 417454
rect 285330 416898 285566 417134
rect 316050 417218 316286 417454
rect 316050 416898 316286 417134
rect 346770 417218 347006 417454
rect 346770 416898 347006 417134
rect 377490 417218 377726 417454
rect 377490 416898 377726 417134
rect 408210 417218 408446 417454
rect 408210 416898 408446 417134
rect 239250 399218 239486 399454
rect 239250 398898 239486 399134
rect 269970 399218 270206 399454
rect 269970 398898 270206 399134
rect 300690 399218 300926 399454
rect 300690 398898 300926 399134
rect 331410 399218 331646 399454
rect 331410 398898 331646 399134
rect 362130 399218 362366 399454
rect 362130 398898 362366 399134
rect 392850 399218 393086 399454
rect 392850 398898 393086 399134
rect 423570 399218 423806 399454
rect 423570 398898 423806 399134
rect 254610 381218 254846 381454
rect 254610 380898 254846 381134
rect 285330 381218 285566 381454
rect 285330 380898 285566 381134
rect 316050 381218 316286 381454
rect 316050 380898 316286 381134
rect 346770 381218 347006 381454
rect 346770 380898 347006 381134
rect 377490 381218 377726 381454
rect 377490 380898 377726 381134
rect 408210 381218 408446 381454
rect 408210 380898 408446 381134
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 300690 363218 300926 363454
rect 300690 362898 300926 363134
rect 331410 363218 331646 363454
rect 331410 362898 331646 363134
rect 362130 363218 362366 363454
rect 362130 362898 362366 363134
rect 392850 363218 393086 363454
rect 392850 362898 393086 363134
rect 423570 363218 423806 363454
rect 423570 362898 423806 363134
rect 254610 345218 254846 345454
rect 254610 344898 254846 345134
rect 285330 345218 285566 345454
rect 285330 344898 285566 345134
rect 316050 345218 316286 345454
rect 316050 344898 316286 345134
rect 346770 345218 347006 345454
rect 346770 344898 347006 345134
rect 377490 345218 377726 345454
rect 377490 344898 377726 345134
rect 408210 345218 408446 345454
rect 408210 344898 408446 345134
rect 239546 312618 240102 313174
rect 239546 276618 240102 277174
rect 239546 240618 240102 241174
rect 239546 204618 240102 205174
rect 239546 168618 240102 169174
rect 239546 132618 240102 133174
rect 239546 96618 240102 97174
rect 239546 60618 240102 61174
rect 235826 20898 236382 21454
rect 235826 -1862 236382 -1306
rect 239546 24618 240102 25174
rect 239546 -3782 240102 -3226
rect 243266 316338 243822 316894
rect 243266 280338 243822 280894
rect 243266 244338 243822 244894
rect 243266 208338 243822 208894
rect 243266 172338 243822 172894
rect 243266 136338 243822 136894
rect 243266 100338 243822 100894
rect 243266 64338 243822 64894
rect 243266 28338 243822 28894
rect 243266 -5702 243822 -5146
rect 246986 320058 247542 320614
rect 246986 284058 247542 284614
rect 246986 248058 247542 248614
rect 246986 212058 247542 212614
rect 246986 176058 247542 176614
rect 246986 140058 247542 140614
rect 246986 104058 247542 104614
rect 246986 68058 247542 68614
rect 246986 32058 247542 32614
rect 228986 -6662 229542 -6106
rect 253826 326898 254382 327454
rect 253826 290898 254382 291454
rect 253826 254898 254382 255454
rect 253826 218898 254382 219454
rect 253826 182898 254382 183454
rect 253826 146898 254382 147454
rect 253826 110898 254382 111454
rect 253826 74898 254382 75454
rect 253826 38898 254382 39454
rect 253826 2898 254382 3454
rect 253826 -902 254382 -346
rect 257546 330618 258102 331174
rect 257546 294618 258102 295174
rect 257546 258618 258102 259174
rect 257546 222618 258102 223174
rect 257546 186618 258102 187174
rect 257546 150618 258102 151174
rect 257546 114618 258102 115174
rect 257546 78618 258102 79174
rect 257546 42618 258102 43174
rect 257546 6618 258102 7174
rect 257546 -2822 258102 -2266
rect 261266 334338 261822 334894
rect 261266 298338 261822 298894
rect 261266 262338 261822 262894
rect 261266 226338 261822 226894
rect 261266 190338 261822 190894
rect 261266 154338 261822 154894
rect 261266 118338 261822 118894
rect 261266 82338 261822 82894
rect 261266 46338 261822 46894
rect 261266 10338 261822 10894
rect 261266 -4742 261822 -4186
rect 264986 302058 265542 302614
rect 264986 266058 265542 266614
rect 264986 230058 265542 230614
rect 264986 194058 265542 194614
rect 264986 158058 265542 158614
rect 264986 122058 265542 122614
rect 264986 86058 265542 86614
rect 264986 50058 265542 50614
rect 264986 14058 265542 14614
rect 246986 -7622 247542 -7066
rect 271826 308898 272382 309454
rect 271826 272898 272382 273454
rect 271826 236898 272382 237454
rect 271826 200898 272382 201454
rect 271826 164898 272382 165454
rect 271826 128898 272382 129454
rect 271826 92898 272382 93454
rect 271826 56898 272382 57454
rect 271826 20898 272382 21454
rect 271826 -1862 272382 -1306
rect 275546 312618 276102 313174
rect 275546 276618 276102 277174
rect 275546 240618 276102 241174
rect 275546 204618 276102 205174
rect 275546 168618 276102 169174
rect 275546 132618 276102 133174
rect 275546 96618 276102 97174
rect 275546 60618 276102 61174
rect 275546 24618 276102 25174
rect 275546 -3782 276102 -3226
rect 279266 316338 279822 316894
rect 279266 280338 279822 280894
rect 279266 244338 279822 244894
rect 279266 208338 279822 208894
rect 279266 172338 279822 172894
rect 279266 136338 279822 136894
rect 279266 100338 279822 100894
rect 279266 64338 279822 64894
rect 279266 28338 279822 28894
rect 279266 -5702 279822 -5146
rect 282986 320058 283542 320614
rect 282986 284058 283542 284614
rect 282986 248058 283542 248614
rect 282986 212058 283542 212614
rect 282986 176058 283542 176614
rect 282986 140058 283542 140614
rect 282986 104058 283542 104614
rect 282986 68058 283542 68614
rect 282986 32058 283542 32614
rect 264986 -6662 265542 -6106
rect 289826 326898 290382 327454
rect 289826 290898 290382 291454
rect 289826 254898 290382 255454
rect 289826 218898 290382 219454
rect 289826 182898 290382 183454
rect 289826 146898 290382 147454
rect 289826 110898 290382 111454
rect 289826 74898 290382 75454
rect 289826 38898 290382 39454
rect 289826 2898 290382 3454
rect 289826 -902 290382 -346
rect 293546 330618 294102 331174
rect 293546 294618 294102 295174
rect 293546 258618 294102 259174
rect 293546 222618 294102 223174
rect 293546 186618 294102 187174
rect 293546 150618 294102 151174
rect 293546 114618 294102 115174
rect 293546 78618 294102 79174
rect 293546 42618 294102 43174
rect 293546 6618 294102 7174
rect 293546 -2822 294102 -2266
rect 297266 334338 297822 334894
rect 297266 298338 297822 298894
rect 297266 262338 297822 262894
rect 297266 226338 297822 226894
rect 297266 190338 297822 190894
rect 297266 154338 297822 154894
rect 297266 118338 297822 118894
rect 297266 82338 297822 82894
rect 297266 46338 297822 46894
rect 297266 10338 297822 10894
rect 297266 -4742 297822 -4186
rect 300986 302058 301542 302614
rect 300986 266058 301542 266614
rect 300986 230058 301542 230614
rect 300986 194058 301542 194614
rect 300986 158058 301542 158614
rect 300986 122058 301542 122614
rect 300986 86058 301542 86614
rect 300986 50058 301542 50614
rect 300986 14058 301542 14614
rect 282986 -7622 283542 -7066
rect 307826 308898 308382 309454
rect 307826 272898 308382 273454
rect 307826 236898 308382 237454
rect 307826 200898 308382 201454
rect 307826 164898 308382 165454
rect 307826 128898 308382 129454
rect 307826 92898 308382 93454
rect 307826 56898 308382 57454
rect 307826 20898 308382 21454
rect 307826 -1862 308382 -1306
rect 311546 312618 312102 313174
rect 311546 276618 312102 277174
rect 311546 240618 312102 241174
rect 311546 204618 312102 205174
rect 311546 168618 312102 169174
rect 311546 132618 312102 133174
rect 311546 96618 312102 97174
rect 311546 60618 312102 61174
rect 311546 24618 312102 25174
rect 311546 -3782 312102 -3226
rect 315266 316338 315822 316894
rect 315266 280338 315822 280894
rect 315266 244338 315822 244894
rect 315266 208338 315822 208894
rect 315266 172338 315822 172894
rect 315266 136338 315822 136894
rect 315266 100338 315822 100894
rect 315266 64338 315822 64894
rect 315266 28338 315822 28894
rect 315266 -5702 315822 -5146
rect 318986 320058 319542 320614
rect 318986 284058 319542 284614
rect 318986 248058 319542 248614
rect 318986 212058 319542 212614
rect 318986 176058 319542 176614
rect 318986 140058 319542 140614
rect 318986 104058 319542 104614
rect 318986 68058 319542 68614
rect 318986 32058 319542 32614
rect 300986 -6662 301542 -6106
rect 325826 326898 326382 327454
rect 325826 290898 326382 291454
rect 325826 254898 326382 255454
rect 325826 218898 326382 219454
rect 325826 182898 326382 183454
rect 325826 146898 326382 147454
rect 325826 110898 326382 111454
rect 325826 74898 326382 75454
rect 325826 38898 326382 39454
rect 325826 2898 326382 3454
rect 325826 -902 326382 -346
rect 329546 330618 330102 331174
rect 329546 294618 330102 295174
rect 329546 258618 330102 259174
rect 329546 222618 330102 223174
rect 329546 186618 330102 187174
rect 329546 150618 330102 151174
rect 329546 114618 330102 115174
rect 329546 78618 330102 79174
rect 329546 42618 330102 43174
rect 329546 6618 330102 7174
rect 329546 -2822 330102 -2266
rect 333266 334338 333822 334894
rect 333266 298338 333822 298894
rect 333266 262338 333822 262894
rect 333266 226338 333822 226894
rect 333266 190338 333822 190894
rect 333266 154338 333822 154894
rect 333266 118338 333822 118894
rect 333266 82338 333822 82894
rect 333266 46338 333822 46894
rect 333266 10338 333822 10894
rect 333266 -4742 333822 -4186
rect 336986 302058 337542 302614
rect 336986 266058 337542 266614
rect 336986 230058 337542 230614
rect 336986 194058 337542 194614
rect 336986 158058 337542 158614
rect 336986 122058 337542 122614
rect 336986 86058 337542 86614
rect 336986 50058 337542 50614
rect 336986 14058 337542 14614
rect 318986 -7622 319542 -7066
rect 343826 308898 344382 309454
rect 343826 272898 344382 273454
rect 343826 236898 344382 237454
rect 343826 200898 344382 201454
rect 343826 164898 344382 165454
rect 343826 128898 344382 129454
rect 343826 92898 344382 93454
rect 343826 56898 344382 57454
rect 343826 20898 344382 21454
rect 343826 -1862 344382 -1306
rect 347546 312618 348102 313174
rect 347546 276618 348102 277174
rect 347546 240618 348102 241174
rect 347546 204618 348102 205174
rect 347546 168618 348102 169174
rect 347546 132618 348102 133174
rect 347546 96618 348102 97174
rect 347546 60618 348102 61174
rect 347546 24618 348102 25174
rect 347546 -3782 348102 -3226
rect 351266 316338 351822 316894
rect 351266 280338 351822 280894
rect 351266 244338 351822 244894
rect 351266 208338 351822 208894
rect 351266 172338 351822 172894
rect 351266 136338 351822 136894
rect 351266 100338 351822 100894
rect 351266 64338 351822 64894
rect 351266 28338 351822 28894
rect 351266 -5702 351822 -5146
rect 354986 320058 355542 320614
rect 354986 284058 355542 284614
rect 354986 248058 355542 248614
rect 354986 212058 355542 212614
rect 354986 176058 355542 176614
rect 354986 140058 355542 140614
rect 354986 104058 355542 104614
rect 354986 68058 355542 68614
rect 354986 32058 355542 32614
rect 336986 -6662 337542 -6106
rect 361826 326898 362382 327454
rect 361826 290898 362382 291454
rect 361826 254898 362382 255454
rect 361826 218898 362382 219454
rect 361826 182898 362382 183454
rect 361826 146898 362382 147454
rect 361826 110898 362382 111454
rect 361826 74898 362382 75454
rect 361826 38898 362382 39454
rect 361826 2898 362382 3454
rect 361826 -902 362382 -346
rect 365546 330618 366102 331174
rect 365546 294618 366102 295174
rect 365546 258618 366102 259174
rect 365546 222618 366102 223174
rect 365546 186618 366102 187174
rect 365546 150618 366102 151174
rect 365546 114618 366102 115174
rect 365546 78618 366102 79174
rect 365546 42618 366102 43174
rect 365546 6618 366102 7174
rect 365546 -2822 366102 -2266
rect 369266 334338 369822 334894
rect 369266 298338 369822 298894
rect 369266 262338 369822 262894
rect 369266 226338 369822 226894
rect 369266 190338 369822 190894
rect 369266 154338 369822 154894
rect 369266 118338 369822 118894
rect 369266 82338 369822 82894
rect 369266 46338 369822 46894
rect 369266 10338 369822 10894
rect 369266 -4742 369822 -4186
rect 372986 302058 373542 302614
rect 372986 266058 373542 266614
rect 372986 230058 373542 230614
rect 372986 194058 373542 194614
rect 372986 158058 373542 158614
rect 372986 122058 373542 122614
rect 372986 86058 373542 86614
rect 372986 50058 373542 50614
rect 372986 14058 373542 14614
rect 354986 -7622 355542 -7066
rect 379826 308898 380382 309454
rect 379826 272898 380382 273454
rect 379826 236898 380382 237454
rect 379826 200898 380382 201454
rect 379826 164898 380382 165454
rect 379826 128898 380382 129454
rect 379826 92898 380382 93454
rect 379826 56898 380382 57454
rect 379826 20898 380382 21454
rect 379826 -1862 380382 -1306
rect 383546 312618 384102 313174
rect 383546 276618 384102 277174
rect 383546 240618 384102 241174
rect 383546 204618 384102 205174
rect 383546 168618 384102 169174
rect 383546 132618 384102 133174
rect 383546 96618 384102 97174
rect 383546 60618 384102 61174
rect 383546 24618 384102 25174
rect 383546 -3782 384102 -3226
rect 387266 316338 387822 316894
rect 387266 280338 387822 280894
rect 387266 244338 387822 244894
rect 387266 208338 387822 208894
rect 387266 172338 387822 172894
rect 387266 136338 387822 136894
rect 387266 100338 387822 100894
rect 387266 64338 387822 64894
rect 387266 28338 387822 28894
rect 387266 -5702 387822 -5146
rect 390986 320058 391542 320614
rect 390986 284058 391542 284614
rect 390986 248058 391542 248614
rect 390986 212058 391542 212614
rect 390986 176058 391542 176614
rect 390986 140058 391542 140614
rect 390986 104058 391542 104614
rect 390986 68058 391542 68614
rect 390986 32058 391542 32614
rect 372986 -6662 373542 -6106
rect 397826 326898 398382 327454
rect 397826 290898 398382 291454
rect 397826 254898 398382 255454
rect 397826 218898 398382 219454
rect 397826 182898 398382 183454
rect 397826 146898 398382 147454
rect 397826 110898 398382 111454
rect 397826 74898 398382 75454
rect 397826 38898 398382 39454
rect 397826 2898 398382 3454
rect 397826 -902 398382 -346
rect 401546 330618 402102 331174
rect 401546 294618 402102 295174
rect 401546 258618 402102 259174
rect 401546 222618 402102 223174
rect 401546 186618 402102 187174
rect 401546 150618 402102 151174
rect 401546 114618 402102 115174
rect 401546 78618 402102 79174
rect 401546 42618 402102 43174
rect 401546 6618 402102 7174
rect 401546 -2822 402102 -2266
rect 405266 334338 405822 334894
rect 405266 298338 405822 298894
rect 405266 262338 405822 262894
rect 405266 226338 405822 226894
rect 405266 190338 405822 190894
rect 405266 154338 405822 154894
rect 405266 118338 405822 118894
rect 405266 82338 405822 82894
rect 405266 46338 405822 46894
rect 405266 10338 405822 10894
rect 405266 -4742 405822 -4186
rect 408986 302058 409542 302614
rect 408986 266058 409542 266614
rect 408986 230058 409542 230614
rect 408986 194058 409542 194614
rect 408986 158058 409542 158614
rect 408986 122058 409542 122614
rect 408986 86058 409542 86614
rect 408986 50058 409542 50614
rect 408986 14058 409542 14614
rect 390986 -7622 391542 -7066
rect 415826 308898 416382 309454
rect 415826 272898 416382 273454
rect 415826 236898 416382 237454
rect 415826 200898 416382 201454
rect 415826 164898 416382 165454
rect 415826 128898 416382 129454
rect 415826 92898 416382 93454
rect 415826 56898 416382 57454
rect 415826 20898 416382 21454
rect 415826 -1862 416382 -1306
rect 419546 312618 420102 313174
rect 419546 276618 420102 277174
rect 419546 240618 420102 241174
rect 419546 204618 420102 205174
rect 419546 168618 420102 169174
rect 419546 132618 420102 133174
rect 419546 96618 420102 97174
rect 419546 60618 420102 61174
rect 419546 24618 420102 25174
rect 419546 -3782 420102 -3226
rect 423266 316338 423822 316894
rect 423266 280338 423822 280894
rect 423266 244338 423822 244894
rect 423266 208338 423822 208894
rect 423266 172338 423822 172894
rect 423266 136338 423822 136894
rect 423266 100338 423822 100894
rect 423266 64338 423822 64894
rect 426986 320058 427542 320614
rect 426986 284058 427542 284614
rect 426986 248058 427542 248614
rect 426986 212058 427542 212614
rect 426986 176058 427542 176614
rect 426986 140058 427542 140614
rect 426986 104058 427542 104614
rect 426986 68058 427542 68614
rect 423266 28338 423822 28894
rect 423266 -5702 423822 -5146
rect 426986 32058 427542 32614
rect 408986 -6662 409542 -6106
rect 437546 474618 438102 475174
rect 437546 438618 438102 439174
rect 437546 402618 438102 403174
rect 437546 366618 438102 367174
rect 433826 326898 434382 327454
rect 433826 290898 434382 291454
rect 433826 254898 434382 255454
rect 433826 218898 434382 219454
rect 433826 182898 434382 183454
rect 433826 146898 434382 147454
rect 433826 110898 434382 111454
rect 433826 74898 434382 75454
rect 433826 38898 434382 39454
rect 433826 2898 434382 3454
rect 433826 -902 434382 -346
rect 437546 330618 438102 331174
rect 437546 294618 438102 295174
rect 437546 258618 438102 259174
rect 437546 222618 438102 223174
rect 437546 186618 438102 187174
rect 437546 150618 438102 151174
rect 437546 114618 438102 115174
rect 437546 78618 438102 79174
rect 437546 42618 438102 43174
rect 437546 6618 438102 7174
rect 437546 -2822 438102 -2266
rect 441266 694338 441822 694894
rect 441266 658338 441822 658894
rect 441266 622338 441822 622894
rect 441266 586338 441822 586894
rect 441266 550338 441822 550894
rect 441266 514338 441822 514894
rect 441266 478338 441822 478894
rect 441266 442338 441822 442894
rect 441266 406338 441822 406894
rect 441266 370338 441822 370894
rect 441266 334338 441822 334894
rect 441266 298338 441822 298894
rect 441266 262338 441822 262894
rect 441266 226338 441822 226894
rect 441266 190338 441822 190894
rect 441266 154338 441822 154894
rect 441266 118338 441822 118894
rect 441266 82338 441822 82894
rect 441266 46338 441822 46894
rect 441266 10338 441822 10894
rect 441266 -4742 441822 -4186
rect 462986 711002 463542 711558
rect 459266 709082 459822 709638
rect 455546 707162 456102 707718
rect 444986 698058 445542 698614
rect 444986 662058 445542 662614
rect 444986 626058 445542 626614
rect 444986 590058 445542 590614
rect 444986 554058 445542 554614
rect 444986 518058 445542 518614
rect 444986 482058 445542 482614
rect 444986 446058 445542 446614
rect 444986 410058 445542 410614
rect 444986 374058 445542 374614
rect 444986 338058 445542 338614
rect 444986 302058 445542 302614
rect 444986 266058 445542 266614
rect 444986 230058 445542 230614
rect 444986 194058 445542 194614
rect 444986 158058 445542 158614
rect 444986 122058 445542 122614
rect 444986 86058 445542 86614
rect 444986 50058 445542 50614
rect 444986 14058 445542 14614
rect 426986 -7622 427542 -7066
rect 451826 705242 452382 705798
rect 451826 668898 452382 669454
rect 451826 632898 452382 633454
rect 451826 596898 452382 597454
rect 451826 560898 452382 561454
rect 451826 524898 452382 525454
rect 451826 488898 452382 489454
rect 451826 452898 452382 453454
rect 451826 416898 452382 417454
rect 451826 380898 452382 381454
rect 451826 344898 452382 345454
rect 451826 308898 452382 309454
rect 451826 272898 452382 273454
rect 451826 236898 452382 237454
rect 451826 200898 452382 201454
rect 451826 164898 452382 165454
rect 451826 128898 452382 129454
rect 451826 92898 452382 93454
rect 451826 56898 452382 57454
rect 451826 20898 452382 21454
rect 451826 -1862 452382 -1306
rect 455546 672618 456102 673174
rect 455546 636618 456102 637174
rect 455546 600618 456102 601174
rect 455546 564618 456102 565174
rect 455546 528618 456102 529174
rect 455546 492618 456102 493174
rect 455546 456618 456102 457174
rect 455546 420618 456102 421174
rect 455546 384618 456102 385174
rect 455546 348618 456102 349174
rect 455546 312618 456102 313174
rect 455546 276618 456102 277174
rect 455546 240618 456102 241174
rect 455546 204618 456102 205174
rect 455546 168618 456102 169174
rect 455546 132618 456102 133174
rect 455546 96618 456102 97174
rect 455546 60618 456102 61174
rect 455546 24618 456102 25174
rect 455546 -3782 456102 -3226
rect 459266 676338 459822 676894
rect 459266 640338 459822 640894
rect 459266 604338 459822 604894
rect 459266 568338 459822 568894
rect 459266 532338 459822 532894
rect 459266 496338 459822 496894
rect 459266 460338 459822 460894
rect 459266 424338 459822 424894
rect 459266 388338 459822 388894
rect 459266 352338 459822 352894
rect 459266 316338 459822 316894
rect 459266 280338 459822 280894
rect 459266 244338 459822 244894
rect 459266 208338 459822 208894
rect 459266 172338 459822 172894
rect 459266 136338 459822 136894
rect 459266 100338 459822 100894
rect 459266 64338 459822 64894
rect 459266 28338 459822 28894
rect 459266 -5702 459822 -5146
rect 480986 710042 481542 710598
rect 477266 708122 477822 708678
rect 473546 706202 474102 706758
rect 462986 680058 463542 680614
rect 462986 644058 463542 644614
rect 462986 608058 463542 608614
rect 462986 572058 463542 572614
rect 462986 536058 463542 536614
rect 462986 500058 463542 500614
rect 462986 464058 463542 464614
rect 462986 428058 463542 428614
rect 462986 392058 463542 392614
rect 462986 356058 463542 356614
rect 462986 320058 463542 320614
rect 462986 284058 463542 284614
rect 462986 248058 463542 248614
rect 462986 212058 463542 212614
rect 462986 176058 463542 176614
rect 462986 140058 463542 140614
rect 462986 104058 463542 104614
rect 462986 68058 463542 68614
rect 462986 32058 463542 32614
rect 444986 -6662 445542 -6106
rect 469826 704282 470382 704838
rect 469826 686898 470382 687454
rect 469826 650898 470382 651454
rect 469826 614898 470382 615454
rect 469826 578898 470382 579454
rect 469826 542898 470382 543454
rect 469826 506898 470382 507454
rect 469826 470898 470382 471454
rect 469826 434898 470382 435454
rect 469826 398898 470382 399454
rect 469826 362898 470382 363454
rect 469826 326898 470382 327454
rect 469826 290898 470382 291454
rect 469826 254898 470382 255454
rect 469826 218898 470382 219454
rect 469826 182898 470382 183454
rect 469826 146898 470382 147454
rect 469826 110898 470382 111454
rect 469826 74898 470382 75454
rect 469826 38898 470382 39454
rect 469826 2898 470382 3454
rect 469826 -902 470382 -346
rect 473546 690618 474102 691174
rect 473546 654618 474102 655174
rect 473546 618618 474102 619174
rect 473546 582618 474102 583174
rect 473546 546618 474102 547174
rect 473546 510618 474102 511174
rect 473546 474618 474102 475174
rect 473546 438618 474102 439174
rect 473546 402618 474102 403174
rect 473546 366618 474102 367174
rect 473546 330618 474102 331174
rect 473546 294618 474102 295174
rect 473546 258618 474102 259174
rect 473546 222618 474102 223174
rect 473546 186618 474102 187174
rect 473546 150618 474102 151174
rect 473546 114618 474102 115174
rect 473546 78618 474102 79174
rect 473546 42618 474102 43174
rect 473546 6618 474102 7174
rect 473546 -2822 474102 -2266
rect 477266 694338 477822 694894
rect 477266 658338 477822 658894
rect 477266 622338 477822 622894
rect 477266 586338 477822 586894
rect 477266 550338 477822 550894
rect 477266 514338 477822 514894
rect 477266 478338 477822 478894
rect 477266 442338 477822 442894
rect 477266 406338 477822 406894
rect 477266 370338 477822 370894
rect 477266 334338 477822 334894
rect 477266 298338 477822 298894
rect 477266 262338 477822 262894
rect 477266 226338 477822 226894
rect 477266 190338 477822 190894
rect 477266 154338 477822 154894
rect 477266 118338 477822 118894
rect 477266 82338 477822 82894
rect 477266 46338 477822 46894
rect 477266 10338 477822 10894
rect 477266 -4742 477822 -4186
rect 498986 711002 499542 711558
rect 495266 709082 495822 709638
rect 491546 707162 492102 707718
rect 480986 698058 481542 698614
rect 480986 662058 481542 662614
rect 480986 626058 481542 626614
rect 480986 590058 481542 590614
rect 480986 554058 481542 554614
rect 480986 518058 481542 518614
rect 480986 482058 481542 482614
rect 480986 446058 481542 446614
rect 480986 410058 481542 410614
rect 480986 374058 481542 374614
rect 480986 338058 481542 338614
rect 480986 302058 481542 302614
rect 480986 266058 481542 266614
rect 480986 230058 481542 230614
rect 480986 194058 481542 194614
rect 480986 158058 481542 158614
rect 480986 122058 481542 122614
rect 480986 86058 481542 86614
rect 480986 50058 481542 50614
rect 480986 14058 481542 14614
rect 462986 -7622 463542 -7066
rect 487826 705242 488382 705798
rect 487826 668898 488382 669454
rect 487826 632898 488382 633454
rect 487826 596898 488382 597454
rect 487826 560898 488382 561454
rect 487826 524898 488382 525454
rect 487826 488898 488382 489454
rect 487826 452898 488382 453454
rect 487826 416898 488382 417454
rect 487826 380898 488382 381454
rect 487826 344898 488382 345454
rect 487826 308898 488382 309454
rect 487826 272898 488382 273454
rect 487826 236898 488382 237454
rect 487826 200898 488382 201454
rect 487826 164898 488382 165454
rect 487826 128898 488382 129454
rect 487826 92898 488382 93454
rect 487826 56898 488382 57454
rect 487826 20898 488382 21454
rect 487826 -1862 488382 -1306
rect 491546 672618 492102 673174
rect 491546 636618 492102 637174
rect 491546 600618 492102 601174
rect 491546 564618 492102 565174
rect 491546 528618 492102 529174
rect 491546 492618 492102 493174
rect 491546 456618 492102 457174
rect 491546 420618 492102 421174
rect 491546 384618 492102 385174
rect 491546 348618 492102 349174
rect 491546 312618 492102 313174
rect 491546 276618 492102 277174
rect 491546 240618 492102 241174
rect 491546 204618 492102 205174
rect 491546 168618 492102 169174
rect 491546 132618 492102 133174
rect 491546 96618 492102 97174
rect 491546 60618 492102 61174
rect 491546 24618 492102 25174
rect 491546 -3782 492102 -3226
rect 495266 676338 495822 676894
rect 495266 640338 495822 640894
rect 495266 604338 495822 604894
rect 495266 568338 495822 568894
rect 495266 532338 495822 532894
rect 495266 496338 495822 496894
rect 495266 460338 495822 460894
rect 495266 424338 495822 424894
rect 495266 388338 495822 388894
rect 495266 352338 495822 352894
rect 495266 316338 495822 316894
rect 495266 280338 495822 280894
rect 495266 244338 495822 244894
rect 495266 208338 495822 208894
rect 495266 172338 495822 172894
rect 495266 136338 495822 136894
rect 495266 100338 495822 100894
rect 495266 64338 495822 64894
rect 495266 28338 495822 28894
rect 495266 -5702 495822 -5146
rect 516986 710042 517542 710598
rect 513266 708122 513822 708678
rect 509546 706202 510102 706758
rect 498986 680058 499542 680614
rect 498986 644058 499542 644614
rect 498986 608058 499542 608614
rect 498986 572058 499542 572614
rect 498986 536058 499542 536614
rect 498986 500058 499542 500614
rect 498986 464058 499542 464614
rect 498986 428058 499542 428614
rect 498986 392058 499542 392614
rect 498986 356058 499542 356614
rect 498986 320058 499542 320614
rect 498986 284058 499542 284614
rect 498986 248058 499542 248614
rect 498986 212058 499542 212614
rect 498986 176058 499542 176614
rect 498986 140058 499542 140614
rect 498986 104058 499542 104614
rect 498986 68058 499542 68614
rect 498986 32058 499542 32614
rect 480986 -6662 481542 -6106
rect 505826 704282 506382 704838
rect 505826 686898 506382 687454
rect 505826 650898 506382 651454
rect 505826 614898 506382 615454
rect 505826 578898 506382 579454
rect 505826 542898 506382 543454
rect 505826 506898 506382 507454
rect 505826 470898 506382 471454
rect 505826 434898 506382 435454
rect 505826 398898 506382 399454
rect 505826 362898 506382 363454
rect 505826 326898 506382 327454
rect 505826 290898 506382 291454
rect 505826 254898 506382 255454
rect 505826 218898 506382 219454
rect 505826 182898 506382 183454
rect 505826 146898 506382 147454
rect 505826 110898 506382 111454
rect 505826 74898 506382 75454
rect 505826 38898 506382 39454
rect 505826 2898 506382 3454
rect 505826 -902 506382 -346
rect 509546 690618 510102 691174
rect 509546 654618 510102 655174
rect 509546 618618 510102 619174
rect 509546 582618 510102 583174
rect 509546 546618 510102 547174
rect 509546 510618 510102 511174
rect 509546 474618 510102 475174
rect 509546 438618 510102 439174
rect 509546 402618 510102 403174
rect 509546 366618 510102 367174
rect 509546 330618 510102 331174
rect 509546 294618 510102 295174
rect 509546 258618 510102 259174
rect 509546 222618 510102 223174
rect 509546 186618 510102 187174
rect 509546 150618 510102 151174
rect 509546 114618 510102 115174
rect 509546 78618 510102 79174
rect 509546 42618 510102 43174
rect 509546 6618 510102 7174
rect 509546 -2822 510102 -2266
rect 513266 694338 513822 694894
rect 513266 658338 513822 658894
rect 513266 622338 513822 622894
rect 513266 586338 513822 586894
rect 513266 550338 513822 550894
rect 513266 514338 513822 514894
rect 513266 478338 513822 478894
rect 513266 442338 513822 442894
rect 513266 406338 513822 406894
rect 513266 370338 513822 370894
rect 513266 334338 513822 334894
rect 513266 298338 513822 298894
rect 513266 262338 513822 262894
rect 513266 226338 513822 226894
rect 513266 190338 513822 190894
rect 513266 154338 513822 154894
rect 513266 118338 513822 118894
rect 513266 82338 513822 82894
rect 513266 46338 513822 46894
rect 513266 10338 513822 10894
rect 513266 -4742 513822 -4186
rect 534986 711002 535542 711558
rect 531266 709082 531822 709638
rect 527546 707162 528102 707718
rect 516986 698058 517542 698614
rect 516986 662058 517542 662614
rect 516986 626058 517542 626614
rect 516986 590058 517542 590614
rect 516986 554058 517542 554614
rect 516986 518058 517542 518614
rect 516986 482058 517542 482614
rect 516986 446058 517542 446614
rect 516986 410058 517542 410614
rect 516986 374058 517542 374614
rect 516986 338058 517542 338614
rect 516986 302058 517542 302614
rect 516986 266058 517542 266614
rect 516986 230058 517542 230614
rect 516986 194058 517542 194614
rect 516986 158058 517542 158614
rect 516986 122058 517542 122614
rect 516986 86058 517542 86614
rect 516986 50058 517542 50614
rect 516986 14058 517542 14614
rect 498986 -7622 499542 -7066
rect 523826 705242 524382 705798
rect 523826 668898 524382 669454
rect 523826 632898 524382 633454
rect 523826 596898 524382 597454
rect 523826 560898 524382 561454
rect 523826 524898 524382 525454
rect 523826 488898 524382 489454
rect 523826 452898 524382 453454
rect 523826 416898 524382 417454
rect 523826 380898 524382 381454
rect 523826 344898 524382 345454
rect 523826 308898 524382 309454
rect 523826 272898 524382 273454
rect 523826 236898 524382 237454
rect 523826 200898 524382 201454
rect 523826 164898 524382 165454
rect 523826 128898 524382 129454
rect 523826 92898 524382 93454
rect 523826 56898 524382 57454
rect 523826 20898 524382 21454
rect 523826 -1862 524382 -1306
rect 527546 672618 528102 673174
rect 527546 636618 528102 637174
rect 527546 600618 528102 601174
rect 527546 564618 528102 565174
rect 527546 528618 528102 529174
rect 527546 492618 528102 493174
rect 527546 456618 528102 457174
rect 527546 420618 528102 421174
rect 527546 384618 528102 385174
rect 527546 348618 528102 349174
rect 527546 312618 528102 313174
rect 527546 276618 528102 277174
rect 527546 240618 528102 241174
rect 527546 204618 528102 205174
rect 527546 168618 528102 169174
rect 527546 132618 528102 133174
rect 527546 96618 528102 97174
rect 527546 60618 528102 61174
rect 527546 24618 528102 25174
rect 527546 -3782 528102 -3226
rect 531266 676338 531822 676894
rect 531266 640338 531822 640894
rect 531266 604338 531822 604894
rect 531266 568338 531822 568894
rect 531266 532338 531822 532894
rect 531266 496338 531822 496894
rect 531266 460338 531822 460894
rect 531266 424338 531822 424894
rect 531266 388338 531822 388894
rect 531266 352338 531822 352894
rect 531266 316338 531822 316894
rect 531266 280338 531822 280894
rect 531266 244338 531822 244894
rect 531266 208338 531822 208894
rect 531266 172338 531822 172894
rect 531266 136338 531822 136894
rect 531266 100338 531822 100894
rect 531266 64338 531822 64894
rect 531266 28338 531822 28894
rect 531266 -5702 531822 -5146
rect 552986 710042 553542 710598
rect 549266 708122 549822 708678
rect 545546 706202 546102 706758
rect 534986 680058 535542 680614
rect 534986 644058 535542 644614
rect 534986 608058 535542 608614
rect 534986 572058 535542 572614
rect 534986 536058 535542 536614
rect 534986 500058 535542 500614
rect 534986 464058 535542 464614
rect 534986 428058 535542 428614
rect 534986 392058 535542 392614
rect 534986 356058 535542 356614
rect 534986 320058 535542 320614
rect 534986 284058 535542 284614
rect 534986 248058 535542 248614
rect 534986 212058 535542 212614
rect 534986 176058 535542 176614
rect 534986 140058 535542 140614
rect 534986 104058 535542 104614
rect 534986 68058 535542 68614
rect 534986 32058 535542 32614
rect 516986 -6662 517542 -6106
rect 541826 704282 542382 704838
rect 541826 686898 542382 687454
rect 541826 650898 542382 651454
rect 541826 614898 542382 615454
rect 541826 578898 542382 579454
rect 541826 542898 542382 543454
rect 541826 506898 542382 507454
rect 541826 470898 542382 471454
rect 541826 434898 542382 435454
rect 541826 398898 542382 399454
rect 541826 362898 542382 363454
rect 541826 326898 542382 327454
rect 541826 290898 542382 291454
rect 541826 254898 542382 255454
rect 541826 218898 542382 219454
rect 541826 182898 542382 183454
rect 541826 146898 542382 147454
rect 541826 110898 542382 111454
rect 541826 74898 542382 75454
rect 541826 38898 542382 39454
rect 541826 2898 542382 3454
rect 541826 -902 542382 -346
rect 545546 690618 546102 691174
rect 545546 654618 546102 655174
rect 545546 618618 546102 619174
rect 545546 582618 546102 583174
rect 545546 546618 546102 547174
rect 545546 510618 546102 511174
rect 545546 474618 546102 475174
rect 545546 438618 546102 439174
rect 545546 402618 546102 403174
rect 545546 366618 546102 367174
rect 545546 330618 546102 331174
rect 545546 294618 546102 295174
rect 545546 258618 546102 259174
rect 545546 222618 546102 223174
rect 545546 186618 546102 187174
rect 545546 150618 546102 151174
rect 545546 114618 546102 115174
rect 545546 78618 546102 79174
rect 545546 42618 546102 43174
rect 545546 6618 546102 7174
rect 545546 -2822 546102 -2266
rect 549266 694338 549822 694894
rect 549266 658338 549822 658894
rect 549266 622338 549822 622894
rect 549266 586338 549822 586894
rect 549266 550338 549822 550894
rect 549266 514338 549822 514894
rect 549266 478338 549822 478894
rect 549266 442338 549822 442894
rect 549266 406338 549822 406894
rect 549266 370338 549822 370894
rect 549266 334338 549822 334894
rect 549266 298338 549822 298894
rect 549266 262338 549822 262894
rect 549266 226338 549822 226894
rect 549266 190338 549822 190894
rect 549266 154338 549822 154894
rect 549266 118338 549822 118894
rect 549266 82338 549822 82894
rect 549266 46338 549822 46894
rect 549266 10338 549822 10894
rect 549266 -4742 549822 -4186
rect 570986 711002 571542 711558
rect 567266 709082 567822 709638
rect 563546 707162 564102 707718
rect 552986 698058 553542 698614
rect 552986 662058 553542 662614
rect 552986 626058 553542 626614
rect 552986 590058 553542 590614
rect 552986 554058 553542 554614
rect 552986 518058 553542 518614
rect 552986 482058 553542 482614
rect 552986 446058 553542 446614
rect 552986 410058 553542 410614
rect 552986 374058 553542 374614
rect 552986 338058 553542 338614
rect 552986 302058 553542 302614
rect 552986 266058 553542 266614
rect 552986 230058 553542 230614
rect 552986 194058 553542 194614
rect 552986 158058 553542 158614
rect 552986 122058 553542 122614
rect 552986 86058 553542 86614
rect 552986 50058 553542 50614
rect 552986 14058 553542 14614
rect 534986 -7622 535542 -7066
rect 559826 705242 560382 705798
rect 559826 668898 560382 669454
rect 559826 632898 560382 633454
rect 559826 596898 560382 597454
rect 559826 560898 560382 561454
rect 559826 524898 560382 525454
rect 559826 488898 560382 489454
rect 559826 452898 560382 453454
rect 559826 416898 560382 417454
rect 559826 380898 560382 381454
rect 559826 344898 560382 345454
rect 559826 308898 560382 309454
rect 559826 272898 560382 273454
rect 559826 236898 560382 237454
rect 559826 200898 560382 201454
rect 559826 164898 560382 165454
rect 559826 128898 560382 129454
rect 559826 92898 560382 93454
rect 559826 56898 560382 57454
rect 559826 20898 560382 21454
rect 559826 -1862 560382 -1306
rect 563546 672618 564102 673174
rect 563546 636618 564102 637174
rect 563546 600618 564102 601174
rect 563546 564618 564102 565174
rect 563546 528618 564102 529174
rect 563546 492618 564102 493174
rect 563546 456618 564102 457174
rect 563546 420618 564102 421174
rect 563546 384618 564102 385174
rect 563546 348618 564102 349174
rect 563546 312618 564102 313174
rect 563546 276618 564102 277174
rect 563546 240618 564102 241174
rect 563546 204618 564102 205174
rect 563546 168618 564102 169174
rect 563546 132618 564102 133174
rect 563546 96618 564102 97174
rect 563546 60618 564102 61174
rect 563546 24618 564102 25174
rect 563546 -3782 564102 -3226
rect 567266 676338 567822 676894
rect 567266 640338 567822 640894
rect 567266 604338 567822 604894
rect 567266 568338 567822 568894
rect 567266 532338 567822 532894
rect 567266 496338 567822 496894
rect 567266 460338 567822 460894
rect 567266 424338 567822 424894
rect 567266 388338 567822 388894
rect 567266 352338 567822 352894
rect 567266 316338 567822 316894
rect 567266 280338 567822 280894
rect 567266 244338 567822 244894
rect 567266 208338 567822 208894
rect 567266 172338 567822 172894
rect 567266 136338 567822 136894
rect 567266 100338 567822 100894
rect 567266 64338 567822 64894
rect 567266 28338 567822 28894
rect 567266 -5702 567822 -5146
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 581546 706202 582102 706758
rect 570986 680058 571542 680614
rect 570986 644058 571542 644614
rect 570986 608058 571542 608614
rect 570986 572058 571542 572614
rect 570986 536058 571542 536614
rect 570986 500058 571542 500614
rect 577826 704282 578382 704838
rect 577826 686898 578382 687454
rect 577826 650898 578382 651454
rect 577826 614898 578382 615454
rect 577826 578898 578382 579454
rect 577826 542898 578382 543454
rect 577826 506898 578382 507454
rect 570986 464058 571542 464614
rect 570986 428058 571542 428614
rect 570986 392058 571542 392614
rect 570986 356058 571542 356614
rect 570986 320058 571542 320614
rect 570986 284058 571542 284614
rect 570986 248058 571542 248614
rect 570986 212058 571542 212614
rect 570986 176058 571542 176614
rect 570986 140058 571542 140614
rect 570986 104058 571542 104614
rect 570986 68058 571542 68614
rect 570986 32058 571542 32614
rect 552986 -6662 553542 -6106
rect 587262 706202 587818 706758
rect 586302 705242 586858 705798
rect 581546 690618 582102 691174
rect 581546 654618 582102 655174
rect 581546 618618 582102 619174
rect 581546 582618 582102 583174
rect 581546 546618 582102 547174
rect 581546 510618 582102 511174
rect 577826 470898 578382 471454
rect 577826 434898 578382 435454
rect 577826 398898 578382 399454
rect 577826 362898 578382 363454
rect 577826 326898 578382 327454
rect 577826 290898 578382 291454
rect 577826 254898 578382 255454
rect 577826 218898 578382 219454
rect 577826 182898 578382 183454
rect 577826 146898 578382 147454
rect 577826 110898 578382 111454
rect 577826 74898 578382 75454
rect 581546 474618 582102 475174
rect 581546 438618 582102 439174
rect 581546 402618 582102 403174
rect 581546 366618 582102 367174
rect 581546 330618 582102 331174
rect 581546 294618 582102 295174
rect 581546 258618 582102 259174
rect 581546 222618 582102 223174
rect 581546 186618 582102 187174
rect 581546 150618 582102 151174
rect 581546 114618 582102 115174
rect 581546 78618 582102 79174
rect 577826 38898 578382 39454
rect 577826 2898 578382 3454
rect 577826 -902 578382 -346
rect 581546 42618 582102 43174
rect 581546 6618 582102 7174
rect 585342 704282 585898 704838
rect 585342 686898 585898 687454
rect 585342 650898 585898 651454
rect 585342 614898 585898 615454
rect 585342 578898 585898 579454
rect 585342 542898 585898 543454
rect 585342 506898 585898 507454
rect 585342 470898 585898 471454
rect 585342 434898 585898 435454
rect 585342 398898 585898 399454
rect 585342 362898 585898 363454
rect 585342 326898 585898 327454
rect 585342 290898 585898 291454
rect 585342 254898 585898 255454
rect 585342 218898 585898 219454
rect 585342 182898 585898 183454
rect 585342 146898 585898 147454
rect 585342 110898 585898 111454
rect 585342 74898 585898 75454
rect 585342 38898 585898 39454
rect 585342 2898 585898 3454
rect 585342 -902 585898 -346
rect 586302 668898 586858 669454
rect 586302 632898 586858 633454
rect 586302 596898 586858 597454
rect 586302 560898 586858 561454
rect 586302 524898 586858 525454
rect 586302 488898 586858 489454
rect 586302 452898 586858 453454
rect 586302 416898 586858 417454
rect 586302 380898 586858 381454
rect 586302 344898 586858 345454
rect 586302 308898 586858 309454
rect 586302 272898 586858 273454
rect 586302 236898 586858 237454
rect 586302 200898 586858 201454
rect 586302 164898 586858 165454
rect 586302 128898 586858 129454
rect 586302 92898 586858 93454
rect 586302 56898 586858 57454
rect 586302 20898 586858 21454
rect 586302 -1862 586858 -1306
rect 587262 690618 587818 691174
rect 587262 654618 587818 655174
rect 587262 618618 587818 619174
rect 587262 582618 587818 583174
rect 587262 546618 587818 547174
rect 587262 510618 587818 511174
rect 587262 474618 587818 475174
rect 587262 438618 587818 439174
rect 587262 402618 587818 403174
rect 587262 366618 587818 367174
rect 587262 330618 587818 331174
rect 587262 294618 587818 295174
rect 587262 258618 587818 259174
rect 587262 222618 587818 223174
rect 587262 186618 587818 187174
rect 587262 150618 587818 151174
rect 587262 114618 587818 115174
rect 587262 78618 587818 79174
rect 587262 42618 587818 43174
rect 587262 6618 587818 7174
rect 581546 -2822 582102 -2266
rect 587262 -2822 587818 -2266
rect 588222 672618 588778 673174
rect 588222 636618 588778 637174
rect 588222 600618 588778 601174
rect 588222 564618 588778 565174
rect 588222 528618 588778 529174
rect 588222 492618 588778 493174
rect 588222 456618 588778 457174
rect 588222 420618 588778 421174
rect 588222 384618 588778 385174
rect 588222 348618 588778 349174
rect 588222 312618 588778 313174
rect 588222 276618 588778 277174
rect 588222 240618 588778 241174
rect 588222 204618 588778 205174
rect 588222 168618 588778 169174
rect 588222 132618 588778 133174
rect 588222 96618 588778 97174
rect 588222 60618 588778 61174
rect 588222 24618 588778 25174
rect 588222 -3782 588778 -3226
rect 589182 694338 589738 694894
rect 589182 658338 589738 658894
rect 589182 622338 589738 622894
rect 589182 586338 589738 586894
rect 589182 550338 589738 550894
rect 589182 514338 589738 514894
rect 589182 478338 589738 478894
rect 589182 442338 589738 442894
rect 589182 406338 589738 406894
rect 589182 370338 589738 370894
rect 589182 334338 589738 334894
rect 589182 298338 589738 298894
rect 589182 262338 589738 262894
rect 589182 226338 589738 226894
rect 589182 190338 589738 190894
rect 589182 154338 589738 154894
rect 589182 118338 589738 118894
rect 589182 82338 589738 82894
rect 589182 46338 589738 46894
rect 589182 10338 589738 10894
rect 589182 -4742 589738 -4186
rect 590142 676338 590698 676894
rect 590142 640338 590698 640894
rect 590142 604338 590698 604894
rect 590142 568338 590698 568894
rect 590142 532338 590698 532894
rect 590142 496338 590698 496894
rect 590142 460338 590698 460894
rect 590142 424338 590698 424894
rect 590142 388338 590698 388894
rect 590142 352338 590698 352894
rect 590142 316338 590698 316894
rect 590142 280338 590698 280894
rect 590142 244338 590698 244894
rect 590142 208338 590698 208894
rect 590142 172338 590698 172894
rect 590142 136338 590698 136894
rect 590142 100338 590698 100894
rect 590142 64338 590698 64894
rect 590142 28338 590698 28894
rect 590142 -5702 590698 -5146
rect 591102 698058 591658 698614
rect 591102 662058 591658 662614
rect 591102 626058 591658 626614
rect 591102 590058 591658 590614
rect 591102 554058 591658 554614
rect 591102 518058 591658 518614
rect 591102 482058 591658 482614
rect 591102 446058 591658 446614
rect 591102 410058 591658 410614
rect 591102 374058 591658 374614
rect 591102 338058 591658 338614
rect 591102 302058 591658 302614
rect 591102 266058 591658 266614
rect 591102 230058 591658 230614
rect 591102 194058 591658 194614
rect 591102 158058 591658 158614
rect 591102 122058 591658 122614
rect 591102 86058 591658 86614
rect 591102 50058 591658 50614
rect 591102 14058 591658 14614
rect 591102 -6662 591658 -6106
rect 592062 680058 592618 680614
rect 592062 644058 592618 644614
rect 592062 608058 592618 608614
rect 592062 572058 592618 572614
rect 592062 536058 592618 536614
rect 592062 500058 592618 500614
rect 592062 464058 592618 464614
rect 592062 428058 592618 428614
rect 592062 392058 592618 392614
rect 592062 356058 592618 356614
rect 592062 320058 592618 320614
rect 592062 284058 592618 284614
rect 592062 248058 592618 248614
rect 592062 212058 592618 212614
rect 592062 176058 592618 176614
rect 592062 140058 592618 140614
rect 592062 104058 592618 104614
rect 592062 68058 592618 68614
rect 592062 32058 592618 32614
rect 570986 -7622 571542 -7066
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 30986 711558
rect 31542 711002 66986 711558
rect 67542 711002 102986 711558
rect 103542 711002 138986 711558
rect 139542 711002 174986 711558
rect 175542 711002 210986 711558
rect 211542 711002 246986 711558
rect 247542 711002 282986 711558
rect 283542 711002 318986 711558
rect 319542 711002 354986 711558
rect 355542 711002 390986 711558
rect 391542 711002 426986 711558
rect 427542 711002 462986 711558
rect 463542 711002 498986 711558
rect 499542 711002 534986 711558
rect 535542 711002 570986 711558
rect 571542 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 12986 710598
rect 13542 710042 48986 710598
rect 49542 710042 84986 710598
rect 85542 710042 120986 710598
rect 121542 710042 156986 710598
rect 157542 710042 192986 710598
rect 193542 710042 228986 710598
rect 229542 710042 264986 710598
rect 265542 710042 300986 710598
rect 301542 710042 336986 710598
rect 337542 710042 372986 710598
rect 373542 710042 408986 710598
rect 409542 710042 444986 710598
rect 445542 710042 480986 710598
rect 481542 710042 516986 710598
rect 517542 710042 552986 710598
rect 553542 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 27266 709638
rect 27822 709082 63266 709638
rect 63822 709082 99266 709638
rect 99822 709082 135266 709638
rect 135822 709082 171266 709638
rect 171822 709082 207266 709638
rect 207822 709082 243266 709638
rect 243822 709082 279266 709638
rect 279822 709082 315266 709638
rect 315822 709082 351266 709638
rect 351822 709082 387266 709638
rect 387822 709082 423266 709638
rect 423822 709082 459266 709638
rect 459822 709082 495266 709638
rect 495822 709082 531266 709638
rect 531822 709082 567266 709638
rect 567822 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 9266 708678
rect 9822 708122 45266 708678
rect 45822 708122 81266 708678
rect 81822 708122 117266 708678
rect 117822 708122 153266 708678
rect 153822 708122 189266 708678
rect 189822 708122 225266 708678
rect 225822 708122 261266 708678
rect 261822 708122 297266 708678
rect 297822 708122 333266 708678
rect 333822 708122 369266 708678
rect 369822 708122 405266 708678
rect 405822 708122 441266 708678
rect 441822 708122 477266 708678
rect 477822 708122 513266 708678
rect 513822 708122 549266 708678
rect 549822 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 23546 707718
rect 24102 707162 59546 707718
rect 60102 707162 95546 707718
rect 96102 707162 131546 707718
rect 132102 707162 167546 707718
rect 168102 707162 203546 707718
rect 204102 707162 239546 707718
rect 240102 707162 275546 707718
rect 276102 707162 311546 707718
rect 312102 707162 347546 707718
rect 348102 707162 383546 707718
rect 384102 707162 419546 707718
rect 420102 707162 455546 707718
rect 456102 707162 491546 707718
rect 492102 707162 527546 707718
rect 528102 707162 563546 707718
rect 564102 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 5546 706758
rect 6102 706202 41546 706758
rect 42102 706202 77546 706758
rect 78102 706202 113546 706758
rect 114102 706202 149546 706758
rect 150102 706202 185546 706758
rect 186102 706202 221546 706758
rect 222102 706202 257546 706758
rect 258102 706202 293546 706758
rect 294102 706202 329546 706758
rect 330102 706202 365546 706758
rect 366102 706202 401546 706758
rect 402102 706202 437546 706758
rect 438102 706202 473546 706758
rect 474102 706202 509546 706758
rect 510102 706202 545546 706758
rect 546102 706202 581546 706758
rect 582102 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 19826 705798
rect 20382 705242 55826 705798
rect 56382 705242 91826 705798
rect 92382 705242 127826 705798
rect 128382 705242 163826 705798
rect 164382 705242 199826 705798
rect 200382 705242 235826 705798
rect 236382 705242 271826 705798
rect 272382 705242 307826 705798
rect 308382 705242 343826 705798
rect 344382 705242 379826 705798
rect 380382 705242 415826 705798
rect 416382 705242 451826 705798
rect 452382 705242 487826 705798
rect 488382 705242 523826 705798
rect 524382 705242 559826 705798
rect 560382 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1826 704838
rect 2382 704282 37826 704838
rect 38382 704282 73826 704838
rect 74382 704282 109826 704838
rect 110382 704282 145826 704838
rect 146382 704282 181826 704838
rect 182382 704282 217826 704838
rect 218382 704282 253826 704838
rect 254382 704282 289826 704838
rect 290382 704282 325826 704838
rect 326382 704282 361826 704838
rect 362382 704282 397826 704838
rect 398382 704282 433826 704838
rect 434382 704282 469826 704838
rect 470382 704282 505826 704838
rect 506382 704282 541826 704838
rect 542382 704282 577826 704838
rect 578382 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698058 -7734 698614
rect -7178 698058 12986 698614
rect 13542 698058 48986 698614
rect 49542 698058 84986 698614
rect 85542 698058 120986 698614
rect 121542 698058 156986 698614
rect 157542 698058 192986 698614
rect 193542 698058 228986 698614
rect 229542 698058 264986 698614
rect 265542 698058 300986 698614
rect 301542 698058 336986 698614
rect 337542 698058 372986 698614
rect 373542 698058 408986 698614
rect 409542 698058 444986 698614
rect 445542 698058 480986 698614
rect 481542 698058 516986 698614
rect 517542 698058 552986 698614
rect 553542 698058 591102 698614
rect 591658 698058 592650 698614
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694338 -5814 694894
rect -5258 694338 9266 694894
rect 9822 694338 45266 694894
rect 45822 694338 81266 694894
rect 81822 694338 117266 694894
rect 117822 694338 153266 694894
rect 153822 694338 189266 694894
rect 189822 694338 225266 694894
rect 225822 694338 261266 694894
rect 261822 694338 297266 694894
rect 297822 694338 333266 694894
rect 333822 694338 369266 694894
rect 369822 694338 405266 694894
rect 405822 694338 441266 694894
rect 441822 694338 477266 694894
rect 477822 694338 513266 694894
rect 513822 694338 549266 694894
rect 549822 694338 589182 694894
rect 589738 694338 590730 694894
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690618 -3894 691174
rect -3338 690618 5546 691174
rect 6102 690618 41546 691174
rect 42102 690618 77546 691174
rect 78102 690618 113546 691174
rect 114102 690618 149546 691174
rect 150102 690618 185546 691174
rect 186102 690618 221546 691174
rect 222102 690618 257546 691174
rect 258102 690618 293546 691174
rect 294102 690618 329546 691174
rect 330102 690618 365546 691174
rect 366102 690618 401546 691174
rect 402102 690618 437546 691174
rect 438102 690618 473546 691174
rect 474102 690618 509546 691174
rect 510102 690618 545546 691174
rect 546102 690618 581546 691174
rect 582102 690618 587262 691174
rect 587818 690618 588810 691174
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 686898 -1974 687454
rect -1418 686898 1826 687454
rect 2382 686898 37826 687454
rect 38382 686898 73826 687454
rect 74382 686898 109826 687454
rect 110382 686898 145826 687454
rect 146382 686898 181826 687454
rect 182382 686898 217826 687454
rect 218382 686898 253826 687454
rect 254382 686898 289826 687454
rect 290382 686898 325826 687454
rect 326382 686898 361826 687454
rect 362382 686898 397826 687454
rect 398382 686898 433826 687454
rect 434382 686898 469826 687454
rect 470382 686898 505826 687454
rect 506382 686898 541826 687454
rect 542382 686898 577826 687454
rect 578382 686898 585342 687454
rect 585898 686898 586890 687454
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680058 -8694 680614
rect -8138 680058 30986 680614
rect 31542 680058 66986 680614
rect 67542 680058 102986 680614
rect 103542 680058 138986 680614
rect 139542 680058 174986 680614
rect 175542 680058 210986 680614
rect 211542 680058 246986 680614
rect 247542 680058 282986 680614
rect 283542 680058 318986 680614
rect 319542 680058 354986 680614
rect 355542 680058 390986 680614
rect 391542 680058 426986 680614
rect 427542 680058 462986 680614
rect 463542 680058 498986 680614
rect 499542 680058 534986 680614
rect 535542 680058 570986 680614
rect 571542 680058 592062 680614
rect 592618 680058 592650 680614
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676338 -6774 676894
rect -6218 676338 27266 676894
rect 27822 676338 63266 676894
rect 63822 676338 99266 676894
rect 99822 676338 135266 676894
rect 135822 676338 171266 676894
rect 171822 676338 207266 676894
rect 207822 676338 243266 676894
rect 243822 676338 279266 676894
rect 279822 676338 315266 676894
rect 315822 676338 351266 676894
rect 351822 676338 387266 676894
rect 387822 676338 423266 676894
rect 423822 676338 459266 676894
rect 459822 676338 495266 676894
rect 495822 676338 531266 676894
rect 531822 676338 567266 676894
rect 567822 676338 590142 676894
rect 590698 676338 590730 676894
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672618 -4854 673174
rect -4298 672618 23546 673174
rect 24102 672618 59546 673174
rect 60102 672618 95546 673174
rect 96102 672618 131546 673174
rect 132102 672618 167546 673174
rect 168102 672618 203546 673174
rect 204102 672618 239546 673174
rect 240102 672618 275546 673174
rect 276102 672618 311546 673174
rect 312102 672618 347546 673174
rect 348102 672618 383546 673174
rect 384102 672618 419546 673174
rect 420102 672618 455546 673174
rect 456102 672618 491546 673174
rect 492102 672618 527546 673174
rect 528102 672618 563546 673174
rect 564102 672618 588222 673174
rect 588778 672618 588810 673174
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 668898 -2934 669454
rect -2378 668898 19826 669454
rect 20382 668898 55826 669454
rect 56382 668898 91826 669454
rect 92382 668898 127826 669454
rect 128382 668898 163826 669454
rect 164382 668898 199826 669454
rect 200382 668898 235826 669454
rect 236382 668898 271826 669454
rect 272382 668898 307826 669454
rect 308382 668898 343826 669454
rect 344382 668898 379826 669454
rect 380382 668898 415826 669454
rect 416382 668898 451826 669454
rect 452382 668898 487826 669454
rect 488382 668898 523826 669454
rect 524382 668898 559826 669454
rect 560382 668898 586302 669454
rect 586858 668898 586890 669454
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662058 -7734 662614
rect -7178 662058 12986 662614
rect 13542 662058 48986 662614
rect 49542 662058 84986 662614
rect 85542 662058 120986 662614
rect 121542 662058 156986 662614
rect 157542 662058 192986 662614
rect 193542 662058 228986 662614
rect 229542 662058 264986 662614
rect 265542 662058 300986 662614
rect 301542 662058 336986 662614
rect 337542 662058 372986 662614
rect 373542 662058 408986 662614
rect 409542 662058 444986 662614
rect 445542 662058 480986 662614
rect 481542 662058 516986 662614
rect 517542 662058 552986 662614
rect 553542 662058 591102 662614
rect 591658 662058 592650 662614
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658338 -5814 658894
rect -5258 658338 9266 658894
rect 9822 658338 45266 658894
rect 45822 658338 81266 658894
rect 81822 658338 117266 658894
rect 117822 658338 153266 658894
rect 153822 658338 189266 658894
rect 189822 658338 225266 658894
rect 225822 658338 261266 658894
rect 261822 658338 297266 658894
rect 297822 658338 333266 658894
rect 333822 658338 369266 658894
rect 369822 658338 405266 658894
rect 405822 658338 441266 658894
rect 441822 658338 477266 658894
rect 477822 658338 513266 658894
rect 513822 658338 549266 658894
rect 549822 658338 589182 658894
rect 589738 658338 590730 658894
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654618 -3894 655174
rect -3338 654618 5546 655174
rect 6102 654618 41546 655174
rect 42102 654618 77546 655174
rect 78102 654618 113546 655174
rect 114102 654618 149546 655174
rect 150102 654618 185546 655174
rect 186102 654618 221546 655174
rect 222102 654618 257546 655174
rect 258102 654618 293546 655174
rect 294102 654618 329546 655174
rect 330102 654618 365546 655174
rect 366102 654618 401546 655174
rect 402102 654618 437546 655174
rect 438102 654618 473546 655174
rect 474102 654618 509546 655174
rect 510102 654618 545546 655174
rect 546102 654618 581546 655174
rect 582102 654618 587262 655174
rect 587818 654618 588810 655174
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 650898 -1974 651454
rect -1418 650898 1826 651454
rect 2382 650898 37826 651454
rect 38382 650898 73826 651454
rect 74382 650898 109826 651454
rect 110382 650898 145826 651454
rect 146382 650898 181826 651454
rect 182382 650898 217826 651454
rect 218382 650898 253826 651454
rect 254382 650898 289826 651454
rect 290382 650898 325826 651454
rect 326382 650898 361826 651454
rect 362382 650898 397826 651454
rect 398382 650898 433826 651454
rect 434382 650898 469826 651454
rect 470382 650898 505826 651454
rect 506382 650898 541826 651454
rect 542382 650898 577826 651454
rect 578382 650898 585342 651454
rect 585898 650898 586890 651454
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644058 -8694 644614
rect -8138 644058 30986 644614
rect 31542 644058 66986 644614
rect 67542 644058 102986 644614
rect 103542 644058 138986 644614
rect 139542 644058 174986 644614
rect 175542 644058 210986 644614
rect 211542 644058 246986 644614
rect 247542 644058 282986 644614
rect 283542 644058 318986 644614
rect 319542 644058 354986 644614
rect 355542 644058 390986 644614
rect 391542 644058 426986 644614
rect 427542 644058 462986 644614
rect 463542 644058 498986 644614
rect 499542 644058 534986 644614
rect 535542 644058 570986 644614
rect 571542 644058 592062 644614
rect 592618 644058 592650 644614
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640338 -6774 640894
rect -6218 640338 27266 640894
rect 27822 640338 63266 640894
rect 63822 640338 99266 640894
rect 99822 640338 135266 640894
rect 135822 640338 171266 640894
rect 171822 640338 207266 640894
rect 207822 640338 243266 640894
rect 243822 640338 279266 640894
rect 279822 640338 315266 640894
rect 315822 640338 351266 640894
rect 351822 640338 387266 640894
rect 387822 640338 423266 640894
rect 423822 640338 459266 640894
rect 459822 640338 495266 640894
rect 495822 640338 531266 640894
rect 531822 640338 567266 640894
rect 567822 640338 590142 640894
rect 590698 640338 590730 640894
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636618 -4854 637174
rect -4298 636618 23546 637174
rect 24102 636618 59546 637174
rect 60102 636618 95546 637174
rect 96102 636618 131546 637174
rect 132102 636618 167546 637174
rect 168102 636618 203546 637174
rect 204102 636618 239546 637174
rect 240102 636618 275546 637174
rect 276102 636618 311546 637174
rect 312102 636618 347546 637174
rect 348102 636618 383546 637174
rect 384102 636618 419546 637174
rect 420102 636618 455546 637174
rect 456102 636618 491546 637174
rect 492102 636618 527546 637174
rect 528102 636618 563546 637174
rect 564102 636618 588222 637174
rect 588778 636618 588810 637174
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 632898 -2934 633454
rect -2378 632898 19826 633454
rect 20382 632898 55826 633454
rect 56382 632898 91826 633454
rect 92382 632898 127826 633454
rect 128382 632898 163826 633454
rect 164382 632898 199826 633454
rect 200382 632898 235826 633454
rect 236382 632898 271826 633454
rect 272382 632898 307826 633454
rect 308382 632898 343826 633454
rect 344382 632898 379826 633454
rect 380382 632898 415826 633454
rect 416382 632898 451826 633454
rect 452382 632898 487826 633454
rect 488382 632898 523826 633454
rect 524382 632898 559826 633454
rect 560382 632898 586302 633454
rect 586858 632898 586890 633454
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626058 -7734 626614
rect -7178 626058 12986 626614
rect 13542 626058 48986 626614
rect 49542 626058 84986 626614
rect 85542 626058 120986 626614
rect 121542 626058 156986 626614
rect 157542 626058 192986 626614
rect 193542 626058 228986 626614
rect 229542 626058 264986 626614
rect 265542 626058 300986 626614
rect 301542 626058 336986 626614
rect 337542 626058 372986 626614
rect 373542 626058 408986 626614
rect 409542 626058 444986 626614
rect 445542 626058 480986 626614
rect 481542 626058 516986 626614
rect 517542 626058 552986 626614
rect 553542 626058 591102 626614
rect 591658 626058 592650 626614
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622338 -5814 622894
rect -5258 622338 9266 622894
rect 9822 622338 45266 622894
rect 45822 622338 81266 622894
rect 81822 622338 117266 622894
rect 117822 622338 153266 622894
rect 153822 622338 189266 622894
rect 189822 622338 225266 622894
rect 225822 622338 261266 622894
rect 261822 622338 297266 622894
rect 297822 622338 333266 622894
rect 333822 622338 369266 622894
rect 369822 622338 405266 622894
rect 405822 622338 441266 622894
rect 441822 622338 477266 622894
rect 477822 622338 513266 622894
rect 513822 622338 549266 622894
rect 549822 622338 589182 622894
rect 589738 622338 590730 622894
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618618 -3894 619174
rect -3338 618618 5546 619174
rect 6102 618618 41546 619174
rect 42102 618618 77546 619174
rect 78102 618618 113546 619174
rect 114102 618618 149546 619174
rect 150102 618618 185546 619174
rect 186102 618618 221546 619174
rect 222102 618618 257546 619174
rect 258102 618618 293546 619174
rect 294102 618618 329546 619174
rect 330102 618618 365546 619174
rect 366102 618618 401546 619174
rect 402102 618618 437546 619174
rect 438102 618618 473546 619174
rect 474102 618618 509546 619174
rect 510102 618618 545546 619174
rect 546102 618618 581546 619174
rect 582102 618618 587262 619174
rect 587818 618618 588810 619174
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 614898 -1974 615454
rect -1418 614898 1826 615454
rect 2382 614898 37826 615454
rect 38382 614898 73826 615454
rect 74382 614898 109826 615454
rect 110382 614898 145826 615454
rect 146382 614898 181826 615454
rect 182382 614898 217826 615454
rect 218382 614898 253826 615454
rect 254382 614898 289826 615454
rect 290382 614898 325826 615454
rect 326382 614898 361826 615454
rect 362382 614898 397826 615454
rect 398382 614898 433826 615454
rect 434382 614898 469826 615454
rect 470382 614898 505826 615454
rect 506382 614898 541826 615454
rect 542382 614898 577826 615454
rect 578382 614898 585342 615454
rect 585898 614898 586890 615454
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608058 -8694 608614
rect -8138 608058 30986 608614
rect 31542 608058 66986 608614
rect 67542 608058 102986 608614
rect 103542 608058 138986 608614
rect 139542 608058 174986 608614
rect 175542 608058 210986 608614
rect 211542 608058 246986 608614
rect 247542 608058 282986 608614
rect 283542 608058 318986 608614
rect 319542 608058 354986 608614
rect 355542 608058 390986 608614
rect 391542 608058 426986 608614
rect 427542 608058 462986 608614
rect 463542 608058 498986 608614
rect 499542 608058 534986 608614
rect 535542 608058 570986 608614
rect 571542 608058 592062 608614
rect 592618 608058 592650 608614
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604338 -6774 604894
rect -6218 604338 27266 604894
rect 27822 604338 63266 604894
rect 63822 604338 99266 604894
rect 99822 604338 135266 604894
rect 135822 604338 171266 604894
rect 171822 604338 207266 604894
rect 207822 604338 243266 604894
rect 243822 604338 279266 604894
rect 279822 604338 315266 604894
rect 315822 604338 351266 604894
rect 351822 604338 387266 604894
rect 387822 604338 423266 604894
rect 423822 604338 459266 604894
rect 459822 604338 495266 604894
rect 495822 604338 531266 604894
rect 531822 604338 567266 604894
rect 567822 604338 590142 604894
rect 590698 604338 590730 604894
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600618 -4854 601174
rect -4298 600618 23546 601174
rect 24102 600618 59546 601174
rect 60102 600618 95546 601174
rect 96102 600618 131546 601174
rect 132102 600618 167546 601174
rect 168102 600618 203546 601174
rect 204102 600618 239546 601174
rect 240102 600618 275546 601174
rect 276102 600618 311546 601174
rect 312102 600618 347546 601174
rect 348102 600618 383546 601174
rect 384102 600618 419546 601174
rect 420102 600618 455546 601174
rect 456102 600618 491546 601174
rect 492102 600618 527546 601174
rect 528102 600618 563546 601174
rect 564102 600618 588222 601174
rect 588778 600618 588810 601174
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 596898 -2934 597454
rect -2378 596898 19826 597454
rect 20382 596898 55826 597454
rect 56382 596898 91826 597454
rect 92382 596898 127826 597454
rect 128382 596898 163826 597454
rect 164382 596898 199826 597454
rect 200382 596898 235826 597454
rect 236382 596898 271826 597454
rect 272382 596898 307826 597454
rect 308382 596898 343826 597454
rect 344382 596898 379826 597454
rect 380382 596898 415826 597454
rect 416382 596898 451826 597454
rect 452382 596898 487826 597454
rect 488382 596898 523826 597454
rect 524382 596898 559826 597454
rect 560382 596898 586302 597454
rect 586858 596898 586890 597454
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590058 -7734 590614
rect -7178 590058 12986 590614
rect 13542 590058 48986 590614
rect 49542 590058 84986 590614
rect 85542 590058 120986 590614
rect 121542 590058 156986 590614
rect 157542 590058 192986 590614
rect 193542 590058 228986 590614
rect 229542 590058 264986 590614
rect 265542 590058 300986 590614
rect 301542 590058 336986 590614
rect 337542 590058 372986 590614
rect 373542 590058 408986 590614
rect 409542 590058 444986 590614
rect 445542 590058 480986 590614
rect 481542 590058 516986 590614
rect 517542 590058 552986 590614
rect 553542 590058 591102 590614
rect 591658 590058 592650 590614
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586338 -5814 586894
rect -5258 586338 9266 586894
rect 9822 586338 45266 586894
rect 45822 586338 81266 586894
rect 81822 586338 117266 586894
rect 117822 586338 153266 586894
rect 153822 586338 189266 586894
rect 189822 586338 225266 586894
rect 225822 586338 261266 586894
rect 261822 586338 297266 586894
rect 297822 586338 333266 586894
rect 333822 586338 369266 586894
rect 369822 586338 405266 586894
rect 405822 586338 441266 586894
rect 441822 586338 477266 586894
rect 477822 586338 513266 586894
rect 513822 586338 549266 586894
rect 549822 586338 589182 586894
rect 589738 586338 590730 586894
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582618 -3894 583174
rect -3338 582618 5546 583174
rect 6102 582618 41546 583174
rect 42102 582618 77546 583174
rect 78102 582618 113546 583174
rect 114102 582618 149546 583174
rect 150102 582618 185546 583174
rect 186102 582618 221546 583174
rect 222102 582618 257546 583174
rect 258102 582618 293546 583174
rect 294102 582618 329546 583174
rect 330102 582618 365546 583174
rect 366102 582618 401546 583174
rect 402102 582618 437546 583174
rect 438102 582618 473546 583174
rect 474102 582618 509546 583174
rect 510102 582618 545546 583174
rect 546102 582618 581546 583174
rect 582102 582618 587262 583174
rect 587818 582618 588810 583174
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 578898 -1974 579454
rect -1418 578898 1826 579454
rect 2382 578898 37826 579454
rect 38382 578898 73826 579454
rect 74382 578898 109826 579454
rect 110382 578898 145826 579454
rect 146382 578898 181826 579454
rect 182382 578898 217826 579454
rect 218382 578898 253826 579454
rect 254382 578898 289826 579454
rect 290382 578898 325826 579454
rect 326382 578898 361826 579454
rect 362382 578898 397826 579454
rect 398382 578898 433826 579454
rect 434382 578898 469826 579454
rect 470382 578898 505826 579454
rect 506382 578898 541826 579454
rect 542382 578898 577826 579454
rect 578382 578898 585342 579454
rect 585898 578898 586890 579454
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572058 -8694 572614
rect -8138 572058 30986 572614
rect 31542 572058 66986 572614
rect 67542 572058 102986 572614
rect 103542 572058 138986 572614
rect 139542 572058 174986 572614
rect 175542 572058 210986 572614
rect 211542 572058 246986 572614
rect 247542 572058 282986 572614
rect 283542 572058 318986 572614
rect 319542 572058 354986 572614
rect 355542 572058 390986 572614
rect 391542 572058 426986 572614
rect 427542 572058 462986 572614
rect 463542 572058 498986 572614
rect 499542 572058 534986 572614
rect 535542 572058 570986 572614
rect 571542 572058 592062 572614
rect 592618 572058 592650 572614
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568338 -6774 568894
rect -6218 568338 27266 568894
rect 27822 568338 63266 568894
rect 63822 568338 99266 568894
rect 99822 568338 135266 568894
rect 135822 568338 171266 568894
rect 171822 568338 207266 568894
rect 207822 568338 243266 568894
rect 243822 568338 279266 568894
rect 279822 568338 315266 568894
rect 315822 568338 351266 568894
rect 351822 568338 387266 568894
rect 387822 568338 423266 568894
rect 423822 568338 459266 568894
rect 459822 568338 495266 568894
rect 495822 568338 531266 568894
rect 531822 568338 567266 568894
rect 567822 568338 590142 568894
rect 590698 568338 590730 568894
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564618 -4854 565174
rect -4298 564618 23546 565174
rect 24102 564618 59546 565174
rect 60102 564618 95546 565174
rect 96102 564618 131546 565174
rect 132102 564618 167546 565174
rect 168102 564618 203546 565174
rect 204102 564618 239546 565174
rect 240102 564618 275546 565174
rect 276102 564618 311546 565174
rect 312102 564618 347546 565174
rect 348102 564618 383546 565174
rect 384102 564618 419546 565174
rect 420102 564618 455546 565174
rect 456102 564618 491546 565174
rect 492102 564618 527546 565174
rect 528102 564618 563546 565174
rect 564102 564618 588222 565174
rect 588778 564618 588810 565174
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 560898 -2934 561454
rect -2378 560898 19826 561454
rect 20382 560898 55826 561454
rect 56382 560898 91826 561454
rect 92382 560898 127826 561454
rect 128382 560898 163826 561454
rect 164382 560898 199826 561454
rect 200382 560898 235826 561454
rect 236382 560898 271826 561454
rect 272382 560898 307826 561454
rect 308382 560898 343826 561454
rect 344382 560898 379826 561454
rect 380382 560898 415826 561454
rect 416382 560898 451826 561454
rect 452382 560898 487826 561454
rect 488382 560898 523826 561454
rect 524382 560898 559826 561454
rect 560382 560898 586302 561454
rect 586858 560898 586890 561454
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554058 -7734 554614
rect -7178 554058 12986 554614
rect 13542 554058 48986 554614
rect 49542 554058 84986 554614
rect 85542 554058 120986 554614
rect 121542 554058 156986 554614
rect 157542 554058 192986 554614
rect 193542 554058 228986 554614
rect 229542 554058 264986 554614
rect 265542 554058 300986 554614
rect 301542 554058 336986 554614
rect 337542 554058 372986 554614
rect 373542 554058 408986 554614
rect 409542 554058 444986 554614
rect 445542 554058 480986 554614
rect 481542 554058 516986 554614
rect 517542 554058 552986 554614
rect 553542 554058 591102 554614
rect 591658 554058 592650 554614
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550338 -5814 550894
rect -5258 550338 9266 550894
rect 9822 550338 45266 550894
rect 45822 550338 81266 550894
rect 81822 550338 117266 550894
rect 117822 550338 153266 550894
rect 153822 550338 189266 550894
rect 189822 550338 225266 550894
rect 225822 550338 261266 550894
rect 261822 550338 297266 550894
rect 297822 550338 333266 550894
rect 333822 550338 369266 550894
rect 369822 550338 405266 550894
rect 405822 550338 441266 550894
rect 441822 550338 477266 550894
rect 477822 550338 513266 550894
rect 513822 550338 549266 550894
rect 549822 550338 589182 550894
rect 589738 550338 590730 550894
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546618 -3894 547174
rect -3338 546618 5546 547174
rect 6102 546618 41546 547174
rect 42102 546618 77546 547174
rect 78102 546618 113546 547174
rect 114102 546618 149546 547174
rect 150102 546618 185546 547174
rect 186102 546618 221546 547174
rect 222102 546618 257546 547174
rect 258102 546618 293546 547174
rect 294102 546618 329546 547174
rect 330102 546618 365546 547174
rect 366102 546618 401546 547174
rect 402102 546618 437546 547174
rect 438102 546618 473546 547174
rect 474102 546618 509546 547174
rect 510102 546618 545546 547174
rect 546102 546618 581546 547174
rect 582102 546618 587262 547174
rect 587818 546618 588810 547174
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 542898 -1974 543454
rect -1418 542898 1826 543454
rect 2382 542898 37826 543454
rect 38382 542898 73826 543454
rect 74382 542898 109826 543454
rect 110382 542898 145826 543454
rect 146382 542898 181826 543454
rect 182382 542898 217826 543454
rect 218382 542898 253826 543454
rect 254382 542898 289826 543454
rect 290382 542898 325826 543454
rect 326382 542898 361826 543454
rect 362382 542898 397826 543454
rect 398382 542898 433826 543454
rect 434382 542898 469826 543454
rect 470382 542898 505826 543454
rect 506382 542898 541826 543454
rect 542382 542898 577826 543454
rect 578382 542898 585342 543454
rect 585898 542898 586890 543454
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536058 -8694 536614
rect -8138 536058 30986 536614
rect 31542 536058 66986 536614
rect 67542 536058 102986 536614
rect 103542 536058 138986 536614
rect 139542 536058 174986 536614
rect 175542 536058 210986 536614
rect 211542 536058 246986 536614
rect 247542 536058 282986 536614
rect 283542 536058 318986 536614
rect 319542 536058 354986 536614
rect 355542 536058 390986 536614
rect 391542 536058 426986 536614
rect 427542 536058 462986 536614
rect 463542 536058 498986 536614
rect 499542 536058 534986 536614
rect 535542 536058 570986 536614
rect 571542 536058 592062 536614
rect 592618 536058 592650 536614
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532338 -6774 532894
rect -6218 532338 27266 532894
rect 27822 532338 63266 532894
rect 63822 532338 99266 532894
rect 99822 532338 135266 532894
rect 135822 532338 171266 532894
rect 171822 532338 207266 532894
rect 207822 532338 243266 532894
rect 243822 532338 279266 532894
rect 279822 532338 315266 532894
rect 315822 532338 351266 532894
rect 351822 532338 387266 532894
rect 387822 532338 423266 532894
rect 423822 532338 459266 532894
rect 459822 532338 495266 532894
rect 495822 532338 531266 532894
rect 531822 532338 567266 532894
rect 567822 532338 590142 532894
rect 590698 532338 590730 532894
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528618 -4854 529174
rect -4298 528618 23546 529174
rect 24102 528618 59546 529174
rect 60102 528618 95546 529174
rect 96102 528618 131546 529174
rect 132102 528618 167546 529174
rect 168102 528618 203546 529174
rect 204102 528618 239546 529174
rect 240102 528618 275546 529174
rect 276102 528618 311546 529174
rect 312102 528618 347546 529174
rect 348102 528618 383546 529174
rect 384102 528618 419546 529174
rect 420102 528618 455546 529174
rect 456102 528618 491546 529174
rect 492102 528618 527546 529174
rect 528102 528618 563546 529174
rect 564102 528618 588222 529174
rect 588778 528618 588810 529174
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 524898 -2934 525454
rect -2378 524898 19826 525454
rect 20382 524898 55826 525454
rect 56382 524898 91826 525454
rect 92382 524898 127826 525454
rect 128382 524898 163826 525454
rect 164382 524898 199826 525454
rect 200382 524898 235826 525454
rect 236382 524898 271826 525454
rect 272382 524898 307826 525454
rect 308382 524898 343826 525454
rect 344382 524898 379826 525454
rect 380382 524898 415826 525454
rect 416382 524898 451826 525454
rect 452382 524898 487826 525454
rect 488382 524898 523826 525454
rect 524382 524898 559826 525454
rect 560382 524898 586302 525454
rect 586858 524898 586890 525454
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518058 -7734 518614
rect -7178 518058 12986 518614
rect 13542 518058 48986 518614
rect 49542 518058 84986 518614
rect 85542 518058 120986 518614
rect 121542 518058 156986 518614
rect 157542 518058 192986 518614
rect 193542 518058 228986 518614
rect 229542 518058 264986 518614
rect 265542 518058 300986 518614
rect 301542 518058 336986 518614
rect 337542 518058 372986 518614
rect 373542 518058 408986 518614
rect 409542 518058 444986 518614
rect 445542 518058 480986 518614
rect 481542 518058 516986 518614
rect 517542 518058 552986 518614
rect 553542 518058 591102 518614
rect 591658 518058 592650 518614
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514338 -5814 514894
rect -5258 514338 9266 514894
rect 9822 514338 45266 514894
rect 45822 514338 81266 514894
rect 81822 514338 117266 514894
rect 117822 514338 153266 514894
rect 153822 514338 189266 514894
rect 189822 514338 225266 514894
rect 225822 514338 261266 514894
rect 261822 514338 297266 514894
rect 297822 514338 333266 514894
rect 333822 514338 369266 514894
rect 369822 514338 405266 514894
rect 405822 514338 441266 514894
rect 441822 514338 477266 514894
rect 477822 514338 513266 514894
rect 513822 514338 549266 514894
rect 549822 514338 589182 514894
rect 589738 514338 590730 514894
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510618 -3894 511174
rect -3338 510618 5546 511174
rect 6102 510618 41546 511174
rect 42102 510618 77546 511174
rect 78102 510618 113546 511174
rect 114102 510618 149546 511174
rect 150102 510618 185546 511174
rect 186102 510618 221546 511174
rect 222102 510618 257546 511174
rect 258102 510618 293546 511174
rect 294102 510618 329546 511174
rect 330102 510618 365546 511174
rect 366102 510618 401546 511174
rect 402102 510618 437546 511174
rect 438102 510618 473546 511174
rect 474102 510618 509546 511174
rect 510102 510618 545546 511174
rect 546102 510618 581546 511174
rect 582102 510618 587262 511174
rect 587818 510618 588810 511174
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 506898 -1974 507454
rect -1418 506898 1826 507454
rect 2382 506898 37826 507454
rect 38382 506898 73826 507454
rect 74382 506898 109826 507454
rect 110382 506898 145826 507454
rect 146382 506898 181826 507454
rect 182382 506898 217826 507454
rect 218382 506898 253826 507454
rect 254382 506898 289826 507454
rect 290382 506898 325826 507454
rect 326382 506898 361826 507454
rect 362382 506898 397826 507454
rect 398382 506898 433826 507454
rect 434382 506898 469826 507454
rect 470382 506898 505826 507454
rect 506382 506898 541826 507454
rect 542382 506898 577826 507454
rect 578382 506898 585342 507454
rect 585898 506898 586890 507454
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500058 -8694 500614
rect -8138 500058 30986 500614
rect 31542 500058 66986 500614
rect 67542 500058 102986 500614
rect 103542 500058 138986 500614
rect 139542 500058 174986 500614
rect 175542 500058 210986 500614
rect 211542 500058 246986 500614
rect 247542 500058 282986 500614
rect 283542 500058 318986 500614
rect 319542 500058 354986 500614
rect 355542 500058 390986 500614
rect 391542 500058 426986 500614
rect 427542 500058 462986 500614
rect 463542 500058 498986 500614
rect 499542 500058 534986 500614
rect 535542 500058 570986 500614
rect 571542 500058 592062 500614
rect 592618 500058 592650 500614
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496338 -6774 496894
rect -6218 496338 27266 496894
rect 27822 496338 63266 496894
rect 63822 496338 99266 496894
rect 99822 496338 135266 496894
rect 135822 496338 171266 496894
rect 171822 496338 207266 496894
rect 207822 496338 459266 496894
rect 459822 496338 495266 496894
rect 495822 496338 531266 496894
rect 531822 496338 567266 496894
rect 567822 496338 590142 496894
rect 590698 496338 590730 496894
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492618 -4854 493174
rect -4298 492618 23546 493174
rect 24102 492618 59546 493174
rect 60102 492618 95546 493174
rect 96102 492618 131546 493174
rect 132102 492618 167546 493174
rect 168102 492618 203546 493174
rect 204102 492618 455546 493174
rect 456102 492618 491546 493174
rect 492102 492618 527546 493174
rect 528102 492618 563546 493174
rect 564102 492618 588222 493174
rect 588778 492618 588810 493174
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 488898 -2934 489454
rect -2378 488898 19826 489454
rect 20382 488898 55826 489454
rect 56382 488898 91826 489454
rect 92382 488898 127826 489454
rect 128382 488898 163826 489454
rect 164382 488898 199826 489454
rect 200382 489218 254610 489454
rect 254846 489218 285330 489454
rect 285566 489218 316050 489454
rect 316286 489218 346770 489454
rect 347006 489218 377490 489454
rect 377726 489218 408210 489454
rect 408446 489218 451826 489454
rect 200382 489134 451826 489218
rect 200382 488898 254610 489134
rect 254846 488898 285330 489134
rect 285566 488898 316050 489134
rect 316286 488898 346770 489134
rect 347006 488898 377490 489134
rect 377726 488898 408210 489134
rect 408446 488898 451826 489134
rect 452382 488898 487826 489454
rect 488382 488898 523826 489454
rect 524382 488898 559826 489454
rect 560382 488898 586302 489454
rect 586858 488898 586890 489454
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482058 -7734 482614
rect -7178 482058 12986 482614
rect 13542 482058 48986 482614
rect 49542 482058 84986 482614
rect 85542 482058 120986 482614
rect 121542 482058 156986 482614
rect 157542 482058 192986 482614
rect 193542 482058 228986 482614
rect 229542 482058 444986 482614
rect 445542 482058 480986 482614
rect 481542 482058 516986 482614
rect 517542 482058 552986 482614
rect 553542 482058 591102 482614
rect 591658 482058 592650 482614
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478338 -5814 478894
rect -5258 478338 9266 478894
rect 9822 478338 45266 478894
rect 45822 478338 81266 478894
rect 81822 478338 117266 478894
rect 117822 478338 153266 478894
rect 153822 478338 189266 478894
rect 189822 478338 225266 478894
rect 225822 478338 441266 478894
rect 441822 478338 477266 478894
rect 477822 478338 513266 478894
rect 513822 478338 549266 478894
rect 549822 478338 589182 478894
rect 589738 478338 590730 478894
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474618 -3894 475174
rect -3338 474618 5546 475174
rect 6102 474618 41546 475174
rect 42102 474618 77546 475174
rect 78102 474618 113546 475174
rect 114102 474618 149546 475174
rect 150102 474618 185546 475174
rect 186102 474618 221546 475174
rect 222102 474618 437546 475174
rect 438102 474618 473546 475174
rect 474102 474618 509546 475174
rect 510102 474618 545546 475174
rect 546102 474618 581546 475174
rect 582102 474618 587262 475174
rect 587818 474618 588810 475174
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 470898 -1974 471454
rect -1418 470898 1826 471454
rect 2382 470898 37826 471454
rect 38382 470898 73826 471454
rect 74382 470898 109826 471454
rect 110382 470898 145826 471454
rect 146382 470898 181826 471454
rect 182382 470898 217826 471454
rect 218382 471218 239250 471454
rect 239486 471218 269970 471454
rect 270206 471218 300690 471454
rect 300926 471218 331410 471454
rect 331646 471218 362130 471454
rect 362366 471218 392850 471454
rect 393086 471218 423570 471454
rect 423806 471218 469826 471454
rect 218382 471134 469826 471218
rect 218382 470898 239250 471134
rect 239486 470898 269970 471134
rect 270206 470898 300690 471134
rect 300926 470898 331410 471134
rect 331646 470898 362130 471134
rect 362366 470898 392850 471134
rect 393086 470898 423570 471134
rect 423806 470898 469826 471134
rect 470382 470898 505826 471454
rect 506382 470898 541826 471454
rect 542382 470898 577826 471454
rect 578382 470898 585342 471454
rect 585898 470898 586890 471454
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464058 -8694 464614
rect -8138 464058 30986 464614
rect 31542 464058 66986 464614
rect 67542 464058 102986 464614
rect 103542 464058 138986 464614
rect 139542 464058 174986 464614
rect 175542 464058 210986 464614
rect 211542 464058 462986 464614
rect 463542 464058 498986 464614
rect 499542 464058 534986 464614
rect 535542 464058 570986 464614
rect 571542 464058 592062 464614
rect 592618 464058 592650 464614
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460338 -6774 460894
rect -6218 460338 27266 460894
rect 27822 460338 63266 460894
rect 63822 460338 99266 460894
rect 99822 460338 135266 460894
rect 135822 460338 171266 460894
rect 171822 460338 207266 460894
rect 207822 460338 459266 460894
rect 459822 460338 495266 460894
rect 495822 460338 531266 460894
rect 531822 460338 567266 460894
rect 567822 460338 590142 460894
rect 590698 460338 590730 460894
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456618 -4854 457174
rect -4298 456618 23546 457174
rect 24102 456618 59546 457174
rect 60102 456618 95546 457174
rect 96102 456618 131546 457174
rect 132102 456618 167546 457174
rect 168102 456618 203546 457174
rect 204102 456618 455546 457174
rect 456102 456618 491546 457174
rect 492102 456618 527546 457174
rect 528102 456618 563546 457174
rect 564102 456618 588222 457174
rect 588778 456618 588810 457174
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 452898 -2934 453454
rect -2378 452898 19826 453454
rect 20382 452898 55826 453454
rect 56382 452898 91826 453454
rect 92382 452898 127826 453454
rect 128382 452898 163826 453454
rect 164382 452898 199826 453454
rect 200382 453218 254610 453454
rect 254846 453218 285330 453454
rect 285566 453218 316050 453454
rect 316286 453218 346770 453454
rect 347006 453218 377490 453454
rect 377726 453218 408210 453454
rect 408446 453218 451826 453454
rect 200382 453134 451826 453218
rect 200382 452898 254610 453134
rect 254846 452898 285330 453134
rect 285566 452898 316050 453134
rect 316286 452898 346770 453134
rect 347006 452898 377490 453134
rect 377726 452898 408210 453134
rect 408446 452898 451826 453134
rect 452382 452898 487826 453454
rect 488382 452898 523826 453454
rect 524382 452898 559826 453454
rect 560382 452898 586302 453454
rect 586858 452898 586890 453454
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446058 -7734 446614
rect -7178 446058 12986 446614
rect 13542 446058 48986 446614
rect 49542 446058 84986 446614
rect 85542 446058 120986 446614
rect 121542 446058 156986 446614
rect 157542 446058 192986 446614
rect 193542 446058 228986 446614
rect 229542 446058 444986 446614
rect 445542 446058 480986 446614
rect 481542 446058 516986 446614
rect 517542 446058 552986 446614
rect 553542 446058 591102 446614
rect 591658 446058 592650 446614
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442338 -5814 442894
rect -5258 442338 9266 442894
rect 9822 442338 45266 442894
rect 45822 442338 81266 442894
rect 81822 442338 117266 442894
rect 117822 442338 153266 442894
rect 153822 442338 189266 442894
rect 189822 442338 225266 442894
rect 225822 442338 441266 442894
rect 441822 442338 477266 442894
rect 477822 442338 513266 442894
rect 513822 442338 549266 442894
rect 549822 442338 589182 442894
rect 589738 442338 590730 442894
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438618 -3894 439174
rect -3338 438618 5546 439174
rect 6102 438618 41546 439174
rect 42102 438618 77546 439174
rect 78102 438618 113546 439174
rect 114102 438618 149546 439174
rect 150102 438618 185546 439174
rect 186102 438618 221546 439174
rect 222102 438618 437546 439174
rect 438102 438618 473546 439174
rect 474102 438618 509546 439174
rect 510102 438618 545546 439174
rect 546102 438618 581546 439174
rect 582102 438618 587262 439174
rect 587818 438618 588810 439174
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 434898 -1974 435454
rect -1418 434898 1826 435454
rect 2382 434898 37826 435454
rect 38382 434898 73826 435454
rect 74382 434898 109826 435454
rect 110382 434898 145826 435454
rect 146382 434898 181826 435454
rect 182382 434898 217826 435454
rect 218382 435218 239250 435454
rect 239486 435218 269970 435454
rect 270206 435218 300690 435454
rect 300926 435218 331410 435454
rect 331646 435218 362130 435454
rect 362366 435218 392850 435454
rect 393086 435218 423570 435454
rect 423806 435218 469826 435454
rect 218382 435134 469826 435218
rect 218382 434898 239250 435134
rect 239486 434898 269970 435134
rect 270206 434898 300690 435134
rect 300926 434898 331410 435134
rect 331646 434898 362130 435134
rect 362366 434898 392850 435134
rect 393086 434898 423570 435134
rect 423806 434898 469826 435134
rect 470382 434898 505826 435454
rect 506382 434898 541826 435454
rect 542382 434898 577826 435454
rect 578382 434898 585342 435454
rect 585898 434898 586890 435454
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428058 -8694 428614
rect -8138 428058 30986 428614
rect 31542 428058 66986 428614
rect 67542 428058 102986 428614
rect 103542 428058 138986 428614
rect 139542 428058 174986 428614
rect 175542 428058 210986 428614
rect 211542 428058 462986 428614
rect 463542 428058 498986 428614
rect 499542 428058 534986 428614
rect 535542 428058 570986 428614
rect 571542 428058 592062 428614
rect 592618 428058 592650 428614
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424338 -6774 424894
rect -6218 424338 27266 424894
rect 27822 424338 63266 424894
rect 63822 424338 99266 424894
rect 99822 424338 135266 424894
rect 135822 424338 171266 424894
rect 171822 424338 207266 424894
rect 207822 424338 459266 424894
rect 459822 424338 495266 424894
rect 495822 424338 531266 424894
rect 531822 424338 567266 424894
rect 567822 424338 590142 424894
rect 590698 424338 590730 424894
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420618 -4854 421174
rect -4298 420618 23546 421174
rect 24102 420618 59546 421174
rect 60102 420618 95546 421174
rect 96102 420618 131546 421174
rect 132102 420618 167546 421174
rect 168102 420618 203546 421174
rect 204102 420618 455546 421174
rect 456102 420618 491546 421174
rect 492102 420618 527546 421174
rect 528102 420618 563546 421174
rect 564102 420618 588222 421174
rect 588778 420618 588810 421174
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 416898 -2934 417454
rect -2378 416898 19826 417454
rect 20382 416898 55826 417454
rect 56382 416898 91826 417454
rect 92382 416898 127826 417454
rect 128382 416898 163826 417454
rect 164382 416898 199826 417454
rect 200382 417218 254610 417454
rect 254846 417218 285330 417454
rect 285566 417218 316050 417454
rect 316286 417218 346770 417454
rect 347006 417218 377490 417454
rect 377726 417218 408210 417454
rect 408446 417218 451826 417454
rect 200382 417134 451826 417218
rect 200382 416898 254610 417134
rect 254846 416898 285330 417134
rect 285566 416898 316050 417134
rect 316286 416898 346770 417134
rect 347006 416898 377490 417134
rect 377726 416898 408210 417134
rect 408446 416898 451826 417134
rect 452382 416898 487826 417454
rect 488382 416898 523826 417454
rect 524382 416898 559826 417454
rect 560382 416898 586302 417454
rect 586858 416898 586890 417454
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410058 -7734 410614
rect -7178 410058 12986 410614
rect 13542 410058 48986 410614
rect 49542 410058 84986 410614
rect 85542 410058 120986 410614
rect 121542 410058 156986 410614
rect 157542 410058 192986 410614
rect 193542 410058 228986 410614
rect 229542 410058 444986 410614
rect 445542 410058 480986 410614
rect 481542 410058 516986 410614
rect 517542 410058 552986 410614
rect 553542 410058 591102 410614
rect 591658 410058 592650 410614
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406338 -5814 406894
rect -5258 406338 9266 406894
rect 9822 406338 45266 406894
rect 45822 406338 81266 406894
rect 81822 406338 117266 406894
rect 117822 406338 153266 406894
rect 153822 406338 189266 406894
rect 189822 406338 225266 406894
rect 225822 406338 441266 406894
rect 441822 406338 477266 406894
rect 477822 406338 513266 406894
rect 513822 406338 549266 406894
rect 549822 406338 589182 406894
rect 589738 406338 590730 406894
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402618 -3894 403174
rect -3338 402618 5546 403174
rect 6102 402618 41546 403174
rect 42102 402618 77546 403174
rect 78102 402618 113546 403174
rect 114102 402618 149546 403174
rect 150102 402618 185546 403174
rect 186102 402618 221546 403174
rect 222102 402618 437546 403174
rect 438102 402618 473546 403174
rect 474102 402618 509546 403174
rect 510102 402618 545546 403174
rect 546102 402618 581546 403174
rect 582102 402618 587262 403174
rect 587818 402618 588810 403174
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 398898 -1974 399454
rect -1418 398898 1826 399454
rect 2382 398898 37826 399454
rect 38382 398898 73826 399454
rect 74382 398898 109826 399454
rect 110382 398898 145826 399454
rect 146382 398898 181826 399454
rect 182382 398898 217826 399454
rect 218382 399218 239250 399454
rect 239486 399218 269970 399454
rect 270206 399218 300690 399454
rect 300926 399218 331410 399454
rect 331646 399218 362130 399454
rect 362366 399218 392850 399454
rect 393086 399218 423570 399454
rect 423806 399218 469826 399454
rect 218382 399134 469826 399218
rect 218382 398898 239250 399134
rect 239486 398898 269970 399134
rect 270206 398898 300690 399134
rect 300926 398898 331410 399134
rect 331646 398898 362130 399134
rect 362366 398898 392850 399134
rect 393086 398898 423570 399134
rect 423806 398898 469826 399134
rect 470382 398898 505826 399454
rect 506382 398898 541826 399454
rect 542382 398898 577826 399454
rect 578382 398898 585342 399454
rect 585898 398898 586890 399454
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392058 -8694 392614
rect -8138 392058 30986 392614
rect 31542 392058 66986 392614
rect 67542 392058 102986 392614
rect 103542 392058 138986 392614
rect 139542 392058 174986 392614
rect 175542 392058 210986 392614
rect 211542 392058 462986 392614
rect 463542 392058 498986 392614
rect 499542 392058 534986 392614
rect 535542 392058 570986 392614
rect 571542 392058 592062 392614
rect 592618 392058 592650 392614
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388338 -6774 388894
rect -6218 388338 27266 388894
rect 27822 388338 63266 388894
rect 63822 388338 99266 388894
rect 99822 388338 135266 388894
rect 135822 388338 171266 388894
rect 171822 388338 207266 388894
rect 207822 388338 459266 388894
rect 459822 388338 495266 388894
rect 495822 388338 531266 388894
rect 531822 388338 567266 388894
rect 567822 388338 590142 388894
rect 590698 388338 590730 388894
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384618 -4854 385174
rect -4298 384618 23546 385174
rect 24102 384618 59546 385174
rect 60102 384618 95546 385174
rect 96102 384618 131546 385174
rect 132102 384618 167546 385174
rect 168102 384618 203546 385174
rect 204102 384618 455546 385174
rect 456102 384618 491546 385174
rect 492102 384618 527546 385174
rect 528102 384618 563546 385174
rect 564102 384618 588222 385174
rect 588778 384618 588810 385174
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 380898 -2934 381454
rect -2378 380898 19826 381454
rect 20382 380898 55826 381454
rect 56382 380898 91826 381454
rect 92382 380898 127826 381454
rect 128382 380898 163826 381454
rect 164382 380898 199826 381454
rect 200382 381218 254610 381454
rect 254846 381218 285330 381454
rect 285566 381218 316050 381454
rect 316286 381218 346770 381454
rect 347006 381218 377490 381454
rect 377726 381218 408210 381454
rect 408446 381218 451826 381454
rect 200382 381134 451826 381218
rect 200382 380898 254610 381134
rect 254846 380898 285330 381134
rect 285566 380898 316050 381134
rect 316286 380898 346770 381134
rect 347006 380898 377490 381134
rect 377726 380898 408210 381134
rect 408446 380898 451826 381134
rect 452382 380898 487826 381454
rect 488382 380898 523826 381454
rect 524382 380898 559826 381454
rect 560382 380898 586302 381454
rect 586858 380898 586890 381454
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374058 -7734 374614
rect -7178 374058 12986 374614
rect 13542 374058 48986 374614
rect 49542 374058 84986 374614
rect 85542 374058 120986 374614
rect 121542 374058 156986 374614
rect 157542 374058 192986 374614
rect 193542 374058 228986 374614
rect 229542 374058 444986 374614
rect 445542 374058 480986 374614
rect 481542 374058 516986 374614
rect 517542 374058 552986 374614
rect 553542 374058 591102 374614
rect 591658 374058 592650 374614
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370338 -5814 370894
rect -5258 370338 9266 370894
rect 9822 370338 45266 370894
rect 45822 370338 81266 370894
rect 81822 370338 117266 370894
rect 117822 370338 153266 370894
rect 153822 370338 189266 370894
rect 189822 370338 225266 370894
rect 225822 370338 441266 370894
rect 441822 370338 477266 370894
rect 477822 370338 513266 370894
rect 513822 370338 549266 370894
rect 549822 370338 589182 370894
rect 589738 370338 590730 370894
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366618 -3894 367174
rect -3338 366618 5546 367174
rect 6102 366618 41546 367174
rect 42102 366618 77546 367174
rect 78102 366618 113546 367174
rect 114102 366618 149546 367174
rect 150102 366618 185546 367174
rect 186102 366618 221546 367174
rect 222102 366618 437546 367174
rect 438102 366618 473546 367174
rect 474102 366618 509546 367174
rect 510102 366618 545546 367174
rect 546102 366618 581546 367174
rect 582102 366618 587262 367174
rect 587818 366618 588810 367174
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 362898 -1974 363454
rect -1418 362898 1826 363454
rect 2382 362898 37826 363454
rect 38382 362898 73826 363454
rect 74382 362898 109826 363454
rect 110382 362898 145826 363454
rect 146382 362898 181826 363454
rect 182382 362898 217826 363454
rect 218382 363218 239250 363454
rect 239486 363218 269970 363454
rect 270206 363218 300690 363454
rect 300926 363218 331410 363454
rect 331646 363218 362130 363454
rect 362366 363218 392850 363454
rect 393086 363218 423570 363454
rect 423806 363218 469826 363454
rect 218382 363134 469826 363218
rect 218382 362898 239250 363134
rect 239486 362898 269970 363134
rect 270206 362898 300690 363134
rect 300926 362898 331410 363134
rect 331646 362898 362130 363134
rect 362366 362898 392850 363134
rect 393086 362898 423570 363134
rect 423806 362898 469826 363134
rect 470382 362898 505826 363454
rect 506382 362898 541826 363454
rect 542382 362898 577826 363454
rect 578382 362898 585342 363454
rect 585898 362898 586890 363454
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356058 -8694 356614
rect -8138 356058 30986 356614
rect 31542 356058 66986 356614
rect 67542 356058 102986 356614
rect 103542 356058 138986 356614
rect 139542 356058 174986 356614
rect 175542 356058 210986 356614
rect 211542 356058 462986 356614
rect 463542 356058 498986 356614
rect 499542 356058 534986 356614
rect 535542 356058 570986 356614
rect 571542 356058 592062 356614
rect 592618 356058 592650 356614
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352338 -6774 352894
rect -6218 352338 27266 352894
rect 27822 352338 63266 352894
rect 63822 352338 99266 352894
rect 99822 352338 135266 352894
rect 135822 352338 171266 352894
rect 171822 352338 207266 352894
rect 207822 352338 459266 352894
rect 459822 352338 495266 352894
rect 495822 352338 531266 352894
rect 531822 352338 567266 352894
rect 567822 352338 590142 352894
rect 590698 352338 590730 352894
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348618 -4854 349174
rect -4298 348618 23546 349174
rect 24102 348618 59546 349174
rect 60102 348618 95546 349174
rect 96102 348618 131546 349174
rect 132102 348618 167546 349174
rect 168102 348618 203546 349174
rect 204102 348618 455546 349174
rect 456102 348618 491546 349174
rect 492102 348618 527546 349174
rect 528102 348618 563546 349174
rect 564102 348618 588222 349174
rect 588778 348618 588810 349174
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 344898 -2934 345454
rect -2378 344898 19826 345454
rect 20382 344898 55826 345454
rect 56382 344898 91826 345454
rect 92382 344898 127826 345454
rect 128382 344898 163826 345454
rect 164382 344898 199826 345454
rect 200382 345218 254610 345454
rect 254846 345218 285330 345454
rect 285566 345218 316050 345454
rect 316286 345218 346770 345454
rect 347006 345218 377490 345454
rect 377726 345218 408210 345454
rect 408446 345218 451826 345454
rect 200382 345134 451826 345218
rect 200382 344898 254610 345134
rect 254846 344898 285330 345134
rect 285566 344898 316050 345134
rect 316286 344898 346770 345134
rect 347006 344898 377490 345134
rect 377726 344898 408210 345134
rect 408446 344898 451826 345134
rect 452382 344898 487826 345454
rect 488382 344898 523826 345454
rect 524382 344898 559826 345454
rect 560382 344898 586302 345454
rect 586858 344898 586890 345454
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338058 -7734 338614
rect -7178 338058 12986 338614
rect 13542 338058 48986 338614
rect 49542 338058 84986 338614
rect 85542 338058 120986 338614
rect 121542 338058 156986 338614
rect 157542 338058 192986 338614
rect 193542 338058 228986 338614
rect 229542 338058 444986 338614
rect 445542 338058 480986 338614
rect 481542 338058 516986 338614
rect 517542 338058 552986 338614
rect 553542 338058 591102 338614
rect 591658 338058 592650 338614
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334338 -5814 334894
rect -5258 334338 9266 334894
rect 9822 334338 45266 334894
rect 45822 334338 81266 334894
rect 81822 334338 117266 334894
rect 117822 334338 153266 334894
rect 153822 334338 189266 334894
rect 189822 334338 225266 334894
rect 225822 334338 261266 334894
rect 261822 334338 297266 334894
rect 297822 334338 333266 334894
rect 333822 334338 369266 334894
rect 369822 334338 405266 334894
rect 405822 334338 441266 334894
rect 441822 334338 477266 334894
rect 477822 334338 513266 334894
rect 513822 334338 549266 334894
rect 549822 334338 589182 334894
rect 589738 334338 590730 334894
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330618 -3894 331174
rect -3338 330618 5546 331174
rect 6102 330618 41546 331174
rect 42102 330618 77546 331174
rect 78102 330618 113546 331174
rect 114102 330618 149546 331174
rect 150102 330618 185546 331174
rect 186102 330618 221546 331174
rect 222102 330618 257546 331174
rect 258102 330618 293546 331174
rect 294102 330618 329546 331174
rect 330102 330618 365546 331174
rect 366102 330618 401546 331174
rect 402102 330618 437546 331174
rect 438102 330618 473546 331174
rect 474102 330618 509546 331174
rect 510102 330618 545546 331174
rect 546102 330618 581546 331174
rect 582102 330618 587262 331174
rect 587818 330618 588810 331174
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 326898 -1974 327454
rect -1418 326898 1826 327454
rect 2382 326898 37826 327454
rect 38382 326898 73826 327454
rect 74382 326898 109826 327454
rect 110382 326898 145826 327454
rect 146382 326898 181826 327454
rect 182382 326898 217826 327454
rect 218382 326898 253826 327454
rect 254382 326898 289826 327454
rect 290382 326898 325826 327454
rect 326382 326898 361826 327454
rect 362382 326898 397826 327454
rect 398382 326898 433826 327454
rect 434382 326898 469826 327454
rect 470382 326898 505826 327454
rect 506382 326898 541826 327454
rect 542382 326898 577826 327454
rect 578382 326898 585342 327454
rect 585898 326898 586890 327454
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320058 -8694 320614
rect -8138 320058 30986 320614
rect 31542 320058 66986 320614
rect 67542 320058 102986 320614
rect 103542 320058 138986 320614
rect 139542 320058 174986 320614
rect 175542 320058 210986 320614
rect 211542 320058 246986 320614
rect 247542 320058 282986 320614
rect 283542 320058 318986 320614
rect 319542 320058 354986 320614
rect 355542 320058 390986 320614
rect 391542 320058 426986 320614
rect 427542 320058 462986 320614
rect 463542 320058 498986 320614
rect 499542 320058 534986 320614
rect 535542 320058 570986 320614
rect 571542 320058 592062 320614
rect 592618 320058 592650 320614
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316338 -6774 316894
rect -6218 316338 27266 316894
rect 27822 316338 63266 316894
rect 63822 316338 99266 316894
rect 99822 316338 135266 316894
rect 135822 316338 171266 316894
rect 171822 316338 207266 316894
rect 207822 316338 243266 316894
rect 243822 316338 279266 316894
rect 279822 316338 315266 316894
rect 315822 316338 351266 316894
rect 351822 316338 387266 316894
rect 387822 316338 423266 316894
rect 423822 316338 459266 316894
rect 459822 316338 495266 316894
rect 495822 316338 531266 316894
rect 531822 316338 567266 316894
rect 567822 316338 590142 316894
rect 590698 316338 590730 316894
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312618 -4854 313174
rect -4298 312618 23546 313174
rect 24102 312618 59546 313174
rect 60102 312618 95546 313174
rect 96102 312618 131546 313174
rect 132102 312618 167546 313174
rect 168102 312618 203546 313174
rect 204102 312618 239546 313174
rect 240102 312618 275546 313174
rect 276102 312618 311546 313174
rect 312102 312618 347546 313174
rect 348102 312618 383546 313174
rect 384102 312618 419546 313174
rect 420102 312618 455546 313174
rect 456102 312618 491546 313174
rect 492102 312618 527546 313174
rect 528102 312618 563546 313174
rect 564102 312618 588222 313174
rect 588778 312618 588810 313174
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 308898 -2934 309454
rect -2378 308898 19826 309454
rect 20382 308898 55826 309454
rect 56382 308898 91826 309454
rect 92382 308898 127826 309454
rect 128382 308898 163826 309454
rect 164382 308898 199826 309454
rect 200382 308898 235826 309454
rect 236382 308898 271826 309454
rect 272382 308898 307826 309454
rect 308382 308898 343826 309454
rect 344382 308898 379826 309454
rect 380382 308898 415826 309454
rect 416382 308898 451826 309454
rect 452382 308898 487826 309454
rect 488382 308898 523826 309454
rect 524382 308898 559826 309454
rect 560382 308898 586302 309454
rect 586858 308898 586890 309454
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302058 -7734 302614
rect -7178 302058 12986 302614
rect 13542 302058 48986 302614
rect 49542 302058 84986 302614
rect 85542 302058 120986 302614
rect 121542 302058 156986 302614
rect 157542 302058 192986 302614
rect 193542 302058 228986 302614
rect 229542 302058 264986 302614
rect 265542 302058 300986 302614
rect 301542 302058 336986 302614
rect 337542 302058 372986 302614
rect 373542 302058 408986 302614
rect 409542 302058 444986 302614
rect 445542 302058 480986 302614
rect 481542 302058 516986 302614
rect 517542 302058 552986 302614
rect 553542 302058 591102 302614
rect 591658 302058 592650 302614
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298338 -5814 298894
rect -5258 298338 9266 298894
rect 9822 298338 45266 298894
rect 45822 298338 81266 298894
rect 81822 298338 117266 298894
rect 117822 298338 153266 298894
rect 153822 298338 189266 298894
rect 189822 298338 225266 298894
rect 225822 298338 261266 298894
rect 261822 298338 297266 298894
rect 297822 298338 333266 298894
rect 333822 298338 369266 298894
rect 369822 298338 405266 298894
rect 405822 298338 441266 298894
rect 441822 298338 477266 298894
rect 477822 298338 513266 298894
rect 513822 298338 549266 298894
rect 549822 298338 589182 298894
rect 589738 298338 590730 298894
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294618 -3894 295174
rect -3338 294618 5546 295174
rect 6102 294618 41546 295174
rect 42102 294618 77546 295174
rect 78102 294618 113546 295174
rect 114102 294618 149546 295174
rect 150102 294618 185546 295174
rect 186102 294618 221546 295174
rect 222102 294618 257546 295174
rect 258102 294618 293546 295174
rect 294102 294618 329546 295174
rect 330102 294618 365546 295174
rect 366102 294618 401546 295174
rect 402102 294618 437546 295174
rect 438102 294618 473546 295174
rect 474102 294618 509546 295174
rect 510102 294618 545546 295174
rect 546102 294618 581546 295174
rect 582102 294618 587262 295174
rect 587818 294618 588810 295174
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 290898 -1974 291454
rect -1418 290898 1826 291454
rect 2382 290898 37826 291454
rect 38382 290898 73826 291454
rect 74382 290898 109826 291454
rect 110382 290898 145826 291454
rect 146382 290898 181826 291454
rect 182382 290898 217826 291454
rect 218382 290898 253826 291454
rect 254382 290898 289826 291454
rect 290382 290898 325826 291454
rect 326382 290898 361826 291454
rect 362382 290898 397826 291454
rect 398382 290898 433826 291454
rect 434382 290898 469826 291454
rect 470382 290898 505826 291454
rect 506382 290898 541826 291454
rect 542382 290898 577826 291454
rect 578382 290898 585342 291454
rect 585898 290898 586890 291454
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284058 -8694 284614
rect -8138 284058 30986 284614
rect 31542 284058 66986 284614
rect 67542 284058 102986 284614
rect 103542 284058 138986 284614
rect 139542 284058 174986 284614
rect 175542 284058 210986 284614
rect 211542 284058 246986 284614
rect 247542 284058 282986 284614
rect 283542 284058 318986 284614
rect 319542 284058 354986 284614
rect 355542 284058 390986 284614
rect 391542 284058 426986 284614
rect 427542 284058 462986 284614
rect 463542 284058 498986 284614
rect 499542 284058 534986 284614
rect 535542 284058 570986 284614
rect 571542 284058 592062 284614
rect 592618 284058 592650 284614
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280338 -6774 280894
rect -6218 280338 27266 280894
rect 27822 280338 63266 280894
rect 63822 280338 99266 280894
rect 99822 280338 135266 280894
rect 135822 280338 171266 280894
rect 171822 280338 207266 280894
rect 207822 280338 243266 280894
rect 243822 280338 279266 280894
rect 279822 280338 315266 280894
rect 315822 280338 351266 280894
rect 351822 280338 387266 280894
rect 387822 280338 423266 280894
rect 423822 280338 459266 280894
rect 459822 280338 495266 280894
rect 495822 280338 531266 280894
rect 531822 280338 567266 280894
rect 567822 280338 590142 280894
rect 590698 280338 590730 280894
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276618 -4854 277174
rect -4298 276618 23546 277174
rect 24102 276618 59546 277174
rect 60102 276618 95546 277174
rect 96102 276618 131546 277174
rect 132102 276618 167546 277174
rect 168102 276618 203546 277174
rect 204102 276618 239546 277174
rect 240102 276618 275546 277174
rect 276102 276618 311546 277174
rect 312102 276618 347546 277174
rect 348102 276618 383546 277174
rect 384102 276618 419546 277174
rect 420102 276618 455546 277174
rect 456102 276618 491546 277174
rect 492102 276618 527546 277174
rect 528102 276618 563546 277174
rect 564102 276618 588222 277174
rect 588778 276618 588810 277174
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 272898 -2934 273454
rect -2378 272898 19826 273454
rect 20382 272898 55826 273454
rect 56382 272898 91826 273454
rect 92382 272898 127826 273454
rect 128382 272898 163826 273454
rect 164382 272898 199826 273454
rect 200382 272898 235826 273454
rect 236382 272898 271826 273454
rect 272382 272898 307826 273454
rect 308382 272898 343826 273454
rect 344382 272898 379826 273454
rect 380382 272898 415826 273454
rect 416382 272898 451826 273454
rect 452382 272898 487826 273454
rect 488382 272898 523826 273454
rect 524382 272898 559826 273454
rect 560382 272898 586302 273454
rect 586858 272898 586890 273454
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266058 -7734 266614
rect -7178 266058 12986 266614
rect 13542 266058 48986 266614
rect 49542 266058 84986 266614
rect 85542 266058 120986 266614
rect 121542 266058 156986 266614
rect 157542 266058 192986 266614
rect 193542 266058 228986 266614
rect 229542 266058 264986 266614
rect 265542 266058 300986 266614
rect 301542 266058 336986 266614
rect 337542 266058 372986 266614
rect 373542 266058 408986 266614
rect 409542 266058 444986 266614
rect 445542 266058 480986 266614
rect 481542 266058 516986 266614
rect 517542 266058 552986 266614
rect 553542 266058 591102 266614
rect 591658 266058 592650 266614
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262338 -5814 262894
rect -5258 262338 9266 262894
rect 9822 262338 45266 262894
rect 45822 262338 81266 262894
rect 81822 262338 117266 262894
rect 117822 262338 153266 262894
rect 153822 262338 189266 262894
rect 189822 262338 225266 262894
rect 225822 262338 261266 262894
rect 261822 262338 297266 262894
rect 297822 262338 333266 262894
rect 333822 262338 369266 262894
rect 369822 262338 405266 262894
rect 405822 262338 441266 262894
rect 441822 262338 477266 262894
rect 477822 262338 513266 262894
rect 513822 262338 549266 262894
rect 549822 262338 589182 262894
rect 589738 262338 590730 262894
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258618 -3894 259174
rect -3338 258618 5546 259174
rect 6102 258618 41546 259174
rect 42102 258618 77546 259174
rect 78102 258618 113546 259174
rect 114102 258618 149546 259174
rect 150102 258618 185546 259174
rect 186102 258618 221546 259174
rect 222102 258618 257546 259174
rect 258102 258618 293546 259174
rect 294102 258618 329546 259174
rect 330102 258618 365546 259174
rect 366102 258618 401546 259174
rect 402102 258618 437546 259174
rect 438102 258618 473546 259174
rect 474102 258618 509546 259174
rect 510102 258618 545546 259174
rect 546102 258618 581546 259174
rect 582102 258618 587262 259174
rect 587818 258618 588810 259174
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 254898 -1974 255454
rect -1418 254898 1826 255454
rect 2382 254898 37826 255454
rect 38382 254898 73826 255454
rect 74382 254898 109826 255454
rect 110382 254898 145826 255454
rect 146382 254898 181826 255454
rect 182382 254898 217826 255454
rect 218382 254898 253826 255454
rect 254382 254898 289826 255454
rect 290382 254898 325826 255454
rect 326382 254898 361826 255454
rect 362382 254898 397826 255454
rect 398382 254898 433826 255454
rect 434382 254898 469826 255454
rect 470382 254898 505826 255454
rect 506382 254898 541826 255454
rect 542382 254898 577826 255454
rect 578382 254898 585342 255454
rect 585898 254898 586890 255454
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248058 -8694 248614
rect -8138 248058 30986 248614
rect 31542 248058 66986 248614
rect 67542 248058 102986 248614
rect 103542 248058 138986 248614
rect 139542 248058 174986 248614
rect 175542 248058 210986 248614
rect 211542 248058 246986 248614
rect 247542 248058 282986 248614
rect 283542 248058 318986 248614
rect 319542 248058 354986 248614
rect 355542 248058 390986 248614
rect 391542 248058 426986 248614
rect 427542 248058 462986 248614
rect 463542 248058 498986 248614
rect 499542 248058 534986 248614
rect 535542 248058 570986 248614
rect 571542 248058 592062 248614
rect 592618 248058 592650 248614
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244338 -6774 244894
rect -6218 244338 27266 244894
rect 27822 244338 63266 244894
rect 63822 244338 99266 244894
rect 99822 244338 135266 244894
rect 135822 244338 171266 244894
rect 171822 244338 207266 244894
rect 207822 244338 243266 244894
rect 243822 244338 279266 244894
rect 279822 244338 315266 244894
rect 315822 244338 351266 244894
rect 351822 244338 387266 244894
rect 387822 244338 423266 244894
rect 423822 244338 459266 244894
rect 459822 244338 495266 244894
rect 495822 244338 531266 244894
rect 531822 244338 567266 244894
rect 567822 244338 590142 244894
rect 590698 244338 590730 244894
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240618 -4854 241174
rect -4298 240618 23546 241174
rect 24102 240618 59546 241174
rect 60102 240618 95546 241174
rect 96102 240618 131546 241174
rect 132102 240618 167546 241174
rect 168102 240618 203546 241174
rect 204102 240618 239546 241174
rect 240102 240618 275546 241174
rect 276102 240618 311546 241174
rect 312102 240618 347546 241174
rect 348102 240618 383546 241174
rect 384102 240618 419546 241174
rect 420102 240618 455546 241174
rect 456102 240618 491546 241174
rect 492102 240618 527546 241174
rect 528102 240618 563546 241174
rect 564102 240618 588222 241174
rect 588778 240618 588810 241174
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 236898 -2934 237454
rect -2378 236898 19826 237454
rect 20382 236898 55826 237454
rect 56382 236898 91826 237454
rect 92382 236898 127826 237454
rect 128382 236898 163826 237454
rect 164382 236898 199826 237454
rect 200382 236898 235826 237454
rect 236382 236898 271826 237454
rect 272382 236898 307826 237454
rect 308382 236898 343826 237454
rect 344382 236898 379826 237454
rect 380382 236898 415826 237454
rect 416382 236898 451826 237454
rect 452382 236898 487826 237454
rect 488382 236898 523826 237454
rect 524382 236898 559826 237454
rect 560382 236898 586302 237454
rect 586858 236898 586890 237454
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230058 -7734 230614
rect -7178 230058 12986 230614
rect 13542 230058 48986 230614
rect 49542 230058 84986 230614
rect 85542 230058 120986 230614
rect 121542 230058 156986 230614
rect 157542 230058 192986 230614
rect 193542 230058 228986 230614
rect 229542 230058 264986 230614
rect 265542 230058 300986 230614
rect 301542 230058 336986 230614
rect 337542 230058 372986 230614
rect 373542 230058 408986 230614
rect 409542 230058 444986 230614
rect 445542 230058 480986 230614
rect 481542 230058 516986 230614
rect 517542 230058 552986 230614
rect 553542 230058 591102 230614
rect 591658 230058 592650 230614
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226338 -5814 226894
rect -5258 226338 9266 226894
rect 9822 226338 45266 226894
rect 45822 226338 81266 226894
rect 81822 226338 117266 226894
rect 117822 226338 153266 226894
rect 153822 226338 189266 226894
rect 189822 226338 225266 226894
rect 225822 226338 261266 226894
rect 261822 226338 297266 226894
rect 297822 226338 333266 226894
rect 333822 226338 369266 226894
rect 369822 226338 405266 226894
rect 405822 226338 441266 226894
rect 441822 226338 477266 226894
rect 477822 226338 513266 226894
rect 513822 226338 549266 226894
rect 549822 226338 589182 226894
rect 589738 226338 590730 226894
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222618 -3894 223174
rect -3338 222618 5546 223174
rect 6102 222618 41546 223174
rect 42102 222618 77546 223174
rect 78102 222618 113546 223174
rect 114102 222618 149546 223174
rect 150102 222618 185546 223174
rect 186102 222618 221546 223174
rect 222102 222618 257546 223174
rect 258102 222618 293546 223174
rect 294102 222618 329546 223174
rect 330102 222618 365546 223174
rect 366102 222618 401546 223174
rect 402102 222618 437546 223174
rect 438102 222618 473546 223174
rect 474102 222618 509546 223174
rect 510102 222618 545546 223174
rect 546102 222618 581546 223174
rect 582102 222618 587262 223174
rect 587818 222618 588810 223174
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 218898 -1974 219454
rect -1418 218898 1826 219454
rect 2382 218898 37826 219454
rect 38382 218898 73826 219454
rect 74382 218898 109826 219454
rect 110382 218898 145826 219454
rect 146382 218898 181826 219454
rect 182382 218898 217826 219454
rect 218382 218898 253826 219454
rect 254382 218898 289826 219454
rect 290382 218898 325826 219454
rect 326382 218898 361826 219454
rect 362382 218898 397826 219454
rect 398382 218898 433826 219454
rect 434382 218898 469826 219454
rect 470382 218898 505826 219454
rect 506382 218898 541826 219454
rect 542382 218898 577826 219454
rect 578382 218898 585342 219454
rect 585898 218898 586890 219454
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212058 -8694 212614
rect -8138 212058 30986 212614
rect 31542 212058 66986 212614
rect 67542 212058 102986 212614
rect 103542 212058 138986 212614
rect 139542 212058 174986 212614
rect 175542 212058 210986 212614
rect 211542 212058 246986 212614
rect 247542 212058 282986 212614
rect 283542 212058 318986 212614
rect 319542 212058 354986 212614
rect 355542 212058 390986 212614
rect 391542 212058 426986 212614
rect 427542 212058 462986 212614
rect 463542 212058 498986 212614
rect 499542 212058 534986 212614
rect 535542 212058 570986 212614
rect 571542 212058 592062 212614
rect 592618 212058 592650 212614
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208338 -6774 208894
rect -6218 208338 27266 208894
rect 27822 208338 63266 208894
rect 63822 208338 99266 208894
rect 99822 208338 135266 208894
rect 135822 208338 171266 208894
rect 171822 208338 207266 208894
rect 207822 208338 243266 208894
rect 243822 208338 279266 208894
rect 279822 208338 315266 208894
rect 315822 208338 351266 208894
rect 351822 208338 387266 208894
rect 387822 208338 423266 208894
rect 423822 208338 459266 208894
rect 459822 208338 495266 208894
rect 495822 208338 531266 208894
rect 531822 208338 567266 208894
rect 567822 208338 590142 208894
rect 590698 208338 590730 208894
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204618 -4854 205174
rect -4298 204618 23546 205174
rect 24102 204618 59546 205174
rect 60102 204618 95546 205174
rect 96102 204618 131546 205174
rect 132102 204618 167546 205174
rect 168102 204618 203546 205174
rect 204102 204618 239546 205174
rect 240102 204618 275546 205174
rect 276102 204618 311546 205174
rect 312102 204618 347546 205174
rect 348102 204618 383546 205174
rect 384102 204618 419546 205174
rect 420102 204618 455546 205174
rect 456102 204618 491546 205174
rect 492102 204618 527546 205174
rect 528102 204618 563546 205174
rect 564102 204618 588222 205174
rect 588778 204618 588810 205174
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 200898 -2934 201454
rect -2378 200898 19826 201454
rect 20382 200898 55826 201454
rect 56382 200898 91826 201454
rect 92382 200898 127826 201454
rect 128382 200898 163826 201454
rect 164382 200898 199826 201454
rect 200382 200898 235826 201454
rect 236382 200898 271826 201454
rect 272382 200898 307826 201454
rect 308382 200898 343826 201454
rect 344382 200898 379826 201454
rect 380382 200898 415826 201454
rect 416382 200898 451826 201454
rect 452382 200898 487826 201454
rect 488382 200898 523826 201454
rect 524382 200898 559826 201454
rect 560382 200898 586302 201454
rect 586858 200898 586890 201454
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194058 -7734 194614
rect -7178 194058 12986 194614
rect 13542 194058 48986 194614
rect 49542 194058 84986 194614
rect 85542 194058 120986 194614
rect 121542 194058 156986 194614
rect 157542 194058 192986 194614
rect 193542 194058 228986 194614
rect 229542 194058 264986 194614
rect 265542 194058 300986 194614
rect 301542 194058 336986 194614
rect 337542 194058 372986 194614
rect 373542 194058 408986 194614
rect 409542 194058 444986 194614
rect 445542 194058 480986 194614
rect 481542 194058 516986 194614
rect 517542 194058 552986 194614
rect 553542 194058 591102 194614
rect 591658 194058 592650 194614
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190338 -5814 190894
rect -5258 190338 9266 190894
rect 9822 190338 45266 190894
rect 45822 190338 81266 190894
rect 81822 190338 117266 190894
rect 117822 190338 153266 190894
rect 153822 190338 189266 190894
rect 189822 190338 225266 190894
rect 225822 190338 261266 190894
rect 261822 190338 297266 190894
rect 297822 190338 333266 190894
rect 333822 190338 369266 190894
rect 369822 190338 405266 190894
rect 405822 190338 441266 190894
rect 441822 190338 477266 190894
rect 477822 190338 513266 190894
rect 513822 190338 549266 190894
rect 549822 190338 589182 190894
rect 589738 190338 590730 190894
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186618 -3894 187174
rect -3338 186618 5546 187174
rect 6102 186618 41546 187174
rect 42102 186618 77546 187174
rect 78102 186618 113546 187174
rect 114102 186618 149546 187174
rect 150102 186618 185546 187174
rect 186102 186618 221546 187174
rect 222102 186618 257546 187174
rect 258102 186618 293546 187174
rect 294102 186618 329546 187174
rect 330102 186618 365546 187174
rect 366102 186618 401546 187174
rect 402102 186618 437546 187174
rect 438102 186618 473546 187174
rect 474102 186618 509546 187174
rect 510102 186618 545546 187174
rect 546102 186618 581546 187174
rect 582102 186618 587262 187174
rect 587818 186618 588810 187174
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 182898 -1974 183454
rect -1418 182898 1826 183454
rect 2382 182898 37826 183454
rect 38382 182898 73826 183454
rect 74382 182898 109826 183454
rect 110382 182898 145826 183454
rect 146382 182898 181826 183454
rect 182382 182898 217826 183454
rect 218382 182898 253826 183454
rect 254382 182898 289826 183454
rect 290382 182898 325826 183454
rect 326382 182898 361826 183454
rect 362382 182898 397826 183454
rect 398382 182898 433826 183454
rect 434382 182898 469826 183454
rect 470382 182898 505826 183454
rect 506382 182898 541826 183454
rect 542382 182898 577826 183454
rect 578382 182898 585342 183454
rect 585898 182898 586890 183454
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176058 -8694 176614
rect -8138 176058 30986 176614
rect 31542 176058 66986 176614
rect 67542 176058 102986 176614
rect 103542 176058 138986 176614
rect 139542 176058 174986 176614
rect 175542 176058 210986 176614
rect 211542 176058 246986 176614
rect 247542 176058 282986 176614
rect 283542 176058 318986 176614
rect 319542 176058 354986 176614
rect 355542 176058 390986 176614
rect 391542 176058 426986 176614
rect 427542 176058 462986 176614
rect 463542 176058 498986 176614
rect 499542 176058 534986 176614
rect 535542 176058 570986 176614
rect 571542 176058 592062 176614
rect 592618 176058 592650 176614
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172338 -6774 172894
rect -6218 172338 27266 172894
rect 27822 172338 63266 172894
rect 63822 172338 99266 172894
rect 99822 172338 135266 172894
rect 135822 172338 171266 172894
rect 171822 172338 207266 172894
rect 207822 172338 243266 172894
rect 243822 172338 279266 172894
rect 279822 172338 315266 172894
rect 315822 172338 351266 172894
rect 351822 172338 387266 172894
rect 387822 172338 423266 172894
rect 423822 172338 459266 172894
rect 459822 172338 495266 172894
rect 495822 172338 531266 172894
rect 531822 172338 567266 172894
rect 567822 172338 590142 172894
rect 590698 172338 590730 172894
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168618 -4854 169174
rect -4298 168618 23546 169174
rect 24102 168618 59546 169174
rect 60102 168618 95546 169174
rect 96102 168618 131546 169174
rect 132102 168618 167546 169174
rect 168102 168618 203546 169174
rect 204102 168618 239546 169174
rect 240102 168618 275546 169174
rect 276102 168618 311546 169174
rect 312102 168618 347546 169174
rect 348102 168618 383546 169174
rect 384102 168618 419546 169174
rect 420102 168618 455546 169174
rect 456102 168618 491546 169174
rect 492102 168618 527546 169174
rect 528102 168618 563546 169174
rect 564102 168618 588222 169174
rect 588778 168618 588810 169174
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 164898 -2934 165454
rect -2378 164898 19826 165454
rect 20382 164898 55826 165454
rect 56382 164898 91826 165454
rect 92382 164898 127826 165454
rect 128382 164898 163826 165454
rect 164382 164898 199826 165454
rect 200382 164898 235826 165454
rect 236382 164898 271826 165454
rect 272382 164898 307826 165454
rect 308382 164898 343826 165454
rect 344382 164898 379826 165454
rect 380382 164898 415826 165454
rect 416382 164898 451826 165454
rect 452382 164898 487826 165454
rect 488382 164898 523826 165454
rect 524382 164898 559826 165454
rect 560382 164898 586302 165454
rect 586858 164898 586890 165454
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158058 -7734 158614
rect -7178 158058 12986 158614
rect 13542 158058 48986 158614
rect 49542 158058 84986 158614
rect 85542 158058 120986 158614
rect 121542 158058 156986 158614
rect 157542 158058 192986 158614
rect 193542 158058 228986 158614
rect 229542 158058 264986 158614
rect 265542 158058 300986 158614
rect 301542 158058 336986 158614
rect 337542 158058 372986 158614
rect 373542 158058 408986 158614
rect 409542 158058 444986 158614
rect 445542 158058 480986 158614
rect 481542 158058 516986 158614
rect 517542 158058 552986 158614
rect 553542 158058 591102 158614
rect 591658 158058 592650 158614
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154338 -5814 154894
rect -5258 154338 9266 154894
rect 9822 154338 45266 154894
rect 45822 154338 81266 154894
rect 81822 154338 117266 154894
rect 117822 154338 153266 154894
rect 153822 154338 189266 154894
rect 189822 154338 225266 154894
rect 225822 154338 261266 154894
rect 261822 154338 297266 154894
rect 297822 154338 333266 154894
rect 333822 154338 369266 154894
rect 369822 154338 405266 154894
rect 405822 154338 441266 154894
rect 441822 154338 477266 154894
rect 477822 154338 513266 154894
rect 513822 154338 549266 154894
rect 549822 154338 589182 154894
rect 589738 154338 590730 154894
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150618 -3894 151174
rect -3338 150618 5546 151174
rect 6102 150618 41546 151174
rect 42102 150618 77546 151174
rect 78102 150618 113546 151174
rect 114102 150618 149546 151174
rect 150102 150618 185546 151174
rect 186102 150618 221546 151174
rect 222102 150618 257546 151174
rect 258102 150618 293546 151174
rect 294102 150618 329546 151174
rect 330102 150618 365546 151174
rect 366102 150618 401546 151174
rect 402102 150618 437546 151174
rect 438102 150618 473546 151174
rect 474102 150618 509546 151174
rect 510102 150618 545546 151174
rect 546102 150618 581546 151174
rect 582102 150618 587262 151174
rect 587818 150618 588810 151174
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 146898 -1974 147454
rect -1418 146898 1826 147454
rect 2382 146898 37826 147454
rect 38382 146898 73826 147454
rect 74382 146898 109826 147454
rect 110382 146898 145826 147454
rect 146382 146898 181826 147454
rect 182382 146898 217826 147454
rect 218382 146898 253826 147454
rect 254382 146898 289826 147454
rect 290382 146898 325826 147454
rect 326382 146898 361826 147454
rect 362382 146898 397826 147454
rect 398382 146898 433826 147454
rect 434382 146898 469826 147454
rect 470382 146898 505826 147454
rect 506382 146898 541826 147454
rect 542382 146898 577826 147454
rect 578382 146898 585342 147454
rect 585898 146898 586890 147454
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140058 -8694 140614
rect -8138 140058 30986 140614
rect 31542 140058 66986 140614
rect 67542 140058 102986 140614
rect 103542 140058 138986 140614
rect 139542 140058 174986 140614
rect 175542 140058 210986 140614
rect 211542 140058 246986 140614
rect 247542 140058 282986 140614
rect 283542 140058 318986 140614
rect 319542 140058 354986 140614
rect 355542 140058 390986 140614
rect 391542 140058 426986 140614
rect 427542 140058 462986 140614
rect 463542 140058 498986 140614
rect 499542 140058 534986 140614
rect 535542 140058 570986 140614
rect 571542 140058 592062 140614
rect 592618 140058 592650 140614
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136338 -6774 136894
rect -6218 136338 27266 136894
rect 27822 136338 63266 136894
rect 63822 136338 99266 136894
rect 99822 136338 135266 136894
rect 135822 136338 171266 136894
rect 171822 136338 207266 136894
rect 207822 136338 243266 136894
rect 243822 136338 279266 136894
rect 279822 136338 315266 136894
rect 315822 136338 351266 136894
rect 351822 136338 387266 136894
rect 387822 136338 423266 136894
rect 423822 136338 459266 136894
rect 459822 136338 495266 136894
rect 495822 136338 531266 136894
rect 531822 136338 567266 136894
rect 567822 136338 590142 136894
rect 590698 136338 590730 136894
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132618 -4854 133174
rect -4298 132618 23546 133174
rect 24102 132618 59546 133174
rect 60102 132618 95546 133174
rect 96102 132618 131546 133174
rect 132102 132618 167546 133174
rect 168102 132618 203546 133174
rect 204102 132618 239546 133174
rect 240102 132618 275546 133174
rect 276102 132618 311546 133174
rect 312102 132618 347546 133174
rect 348102 132618 383546 133174
rect 384102 132618 419546 133174
rect 420102 132618 455546 133174
rect 456102 132618 491546 133174
rect 492102 132618 527546 133174
rect 528102 132618 563546 133174
rect 564102 132618 588222 133174
rect 588778 132618 588810 133174
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 128898 -2934 129454
rect -2378 128898 19826 129454
rect 20382 128898 55826 129454
rect 56382 128898 91826 129454
rect 92382 128898 127826 129454
rect 128382 128898 163826 129454
rect 164382 128898 199826 129454
rect 200382 128898 235826 129454
rect 236382 128898 271826 129454
rect 272382 128898 307826 129454
rect 308382 128898 343826 129454
rect 344382 128898 379826 129454
rect 380382 128898 415826 129454
rect 416382 128898 451826 129454
rect 452382 128898 487826 129454
rect 488382 128898 523826 129454
rect 524382 128898 559826 129454
rect 560382 128898 586302 129454
rect 586858 128898 586890 129454
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122058 -7734 122614
rect -7178 122058 12986 122614
rect 13542 122058 48986 122614
rect 49542 122058 84986 122614
rect 85542 122058 120986 122614
rect 121542 122058 156986 122614
rect 157542 122058 192986 122614
rect 193542 122058 228986 122614
rect 229542 122058 264986 122614
rect 265542 122058 300986 122614
rect 301542 122058 336986 122614
rect 337542 122058 372986 122614
rect 373542 122058 408986 122614
rect 409542 122058 444986 122614
rect 445542 122058 480986 122614
rect 481542 122058 516986 122614
rect 517542 122058 552986 122614
rect 553542 122058 591102 122614
rect 591658 122058 592650 122614
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118338 -5814 118894
rect -5258 118338 9266 118894
rect 9822 118338 45266 118894
rect 45822 118338 81266 118894
rect 81822 118338 117266 118894
rect 117822 118338 153266 118894
rect 153822 118338 189266 118894
rect 189822 118338 225266 118894
rect 225822 118338 261266 118894
rect 261822 118338 297266 118894
rect 297822 118338 333266 118894
rect 333822 118338 369266 118894
rect 369822 118338 405266 118894
rect 405822 118338 441266 118894
rect 441822 118338 477266 118894
rect 477822 118338 513266 118894
rect 513822 118338 549266 118894
rect 549822 118338 589182 118894
rect 589738 118338 590730 118894
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114618 -3894 115174
rect -3338 114618 5546 115174
rect 6102 114618 41546 115174
rect 42102 114618 77546 115174
rect 78102 114618 113546 115174
rect 114102 114618 149546 115174
rect 150102 114618 185546 115174
rect 186102 114618 221546 115174
rect 222102 114618 257546 115174
rect 258102 114618 293546 115174
rect 294102 114618 329546 115174
rect 330102 114618 365546 115174
rect 366102 114618 401546 115174
rect 402102 114618 437546 115174
rect 438102 114618 473546 115174
rect 474102 114618 509546 115174
rect 510102 114618 545546 115174
rect 546102 114618 581546 115174
rect 582102 114618 587262 115174
rect 587818 114618 588810 115174
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 110898 -1974 111454
rect -1418 110898 1826 111454
rect 2382 110898 37826 111454
rect 38382 110898 73826 111454
rect 74382 110898 109826 111454
rect 110382 110898 145826 111454
rect 146382 110898 181826 111454
rect 182382 110898 217826 111454
rect 218382 110898 253826 111454
rect 254382 110898 289826 111454
rect 290382 110898 325826 111454
rect 326382 110898 361826 111454
rect 362382 110898 397826 111454
rect 398382 110898 433826 111454
rect 434382 110898 469826 111454
rect 470382 110898 505826 111454
rect 506382 110898 541826 111454
rect 542382 110898 577826 111454
rect 578382 110898 585342 111454
rect 585898 110898 586890 111454
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104058 -8694 104614
rect -8138 104058 30986 104614
rect 31542 104058 66986 104614
rect 67542 104058 102986 104614
rect 103542 104058 138986 104614
rect 139542 104058 174986 104614
rect 175542 104058 210986 104614
rect 211542 104058 246986 104614
rect 247542 104058 282986 104614
rect 283542 104058 318986 104614
rect 319542 104058 354986 104614
rect 355542 104058 390986 104614
rect 391542 104058 426986 104614
rect 427542 104058 462986 104614
rect 463542 104058 498986 104614
rect 499542 104058 534986 104614
rect 535542 104058 570986 104614
rect 571542 104058 592062 104614
rect 592618 104058 592650 104614
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100338 -6774 100894
rect -6218 100338 27266 100894
rect 27822 100338 63266 100894
rect 63822 100338 99266 100894
rect 99822 100338 135266 100894
rect 135822 100338 171266 100894
rect 171822 100338 207266 100894
rect 207822 100338 243266 100894
rect 243822 100338 279266 100894
rect 279822 100338 315266 100894
rect 315822 100338 351266 100894
rect 351822 100338 387266 100894
rect 387822 100338 423266 100894
rect 423822 100338 459266 100894
rect 459822 100338 495266 100894
rect 495822 100338 531266 100894
rect 531822 100338 567266 100894
rect 567822 100338 590142 100894
rect 590698 100338 590730 100894
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96618 -4854 97174
rect -4298 96618 23546 97174
rect 24102 96618 59546 97174
rect 60102 96618 95546 97174
rect 96102 96618 131546 97174
rect 132102 96618 167546 97174
rect 168102 96618 203546 97174
rect 204102 96618 239546 97174
rect 240102 96618 275546 97174
rect 276102 96618 311546 97174
rect 312102 96618 347546 97174
rect 348102 96618 383546 97174
rect 384102 96618 419546 97174
rect 420102 96618 455546 97174
rect 456102 96618 491546 97174
rect 492102 96618 527546 97174
rect 528102 96618 563546 97174
rect 564102 96618 588222 97174
rect 588778 96618 588810 97174
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 92898 -2934 93454
rect -2378 92898 19826 93454
rect 20382 92898 55826 93454
rect 56382 92898 91826 93454
rect 92382 92898 127826 93454
rect 128382 92898 163826 93454
rect 164382 92898 199826 93454
rect 200382 92898 235826 93454
rect 236382 92898 271826 93454
rect 272382 92898 307826 93454
rect 308382 92898 343826 93454
rect 344382 92898 379826 93454
rect 380382 92898 415826 93454
rect 416382 92898 451826 93454
rect 452382 92898 487826 93454
rect 488382 92898 523826 93454
rect 524382 92898 559826 93454
rect 560382 92898 586302 93454
rect 586858 92898 586890 93454
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86058 -7734 86614
rect -7178 86058 12986 86614
rect 13542 86058 48986 86614
rect 49542 86058 84986 86614
rect 85542 86058 120986 86614
rect 121542 86058 156986 86614
rect 157542 86058 192986 86614
rect 193542 86058 228986 86614
rect 229542 86058 264986 86614
rect 265542 86058 300986 86614
rect 301542 86058 336986 86614
rect 337542 86058 372986 86614
rect 373542 86058 408986 86614
rect 409542 86058 444986 86614
rect 445542 86058 480986 86614
rect 481542 86058 516986 86614
rect 517542 86058 552986 86614
rect 553542 86058 591102 86614
rect 591658 86058 592650 86614
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82338 -5814 82894
rect -5258 82338 9266 82894
rect 9822 82338 45266 82894
rect 45822 82338 81266 82894
rect 81822 82338 117266 82894
rect 117822 82338 153266 82894
rect 153822 82338 189266 82894
rect 189822 82338 225266 82894
rect 225822 82338 261266 82894
rect 261822 82338 297266 82894
rect 297822 82338 333266 82894
rect 333822 82338 369266 82894
rect 369822 82338 405266 82894
rect 405822 82338 441266 82894
rect 441822 82338 477266 82894
rect 477822 82338 513266 82894
rect 513822 82338 549266 82894
rect 549822 82338 589182 82894
rect 589738 82338 590730 82894
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78618 -3894 79174
rect -3338 78618 5546 79174
rect 6102 78618 41546 79174
rect 42102 78618 77546 79174
rect 78102 78618 113546 79174
rect 114102 78618 149546 79174
rect 150102 78618 185546 79174
rect 186102 78618 221546 79174
rect 222102 78618 257546 79174
rect 258102 78618 293546 79174
rect 294102 78618 329546 79174
rect 330102 78618 365546 79174
rect 366102 78618 401546 79174
rect 402102 78618 437546 79174
rect 438102 78618 473546 79174
rect 474102 78618 509546 79174
rect 510102 78618 545546 79174
rect 546102 78618 581546 79174
rect 582102 78618 587262 79174
rect 587818 78618 588810 79174
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 74898 -1974 75454
rect -1418 74898 1826 75454
rect 2382 74898 37826 75454
rect 38382 74898 73826 75454
rect 74382 74898 109826 75454
rect 110382 74898 145826 75454
rect 146382 74898 181826 75454
rect 182382 74898 217826 75454
rect 218382 74898 253826 75454
rect 254382 74898 289826 75454
rect 290382 74898 325826 75454
rect 326382 74898 361826 75454
rect 362382 74898 397826 75454
rect 398382 74898 433826 75454
rect 434382 74898 469826 75454
rect 470382 74898 505826 75454
rect 506382 74898 541826 75454
rect 542382 74898 577826 75454
rect 578382 74898 585342 75454
rect 585898 74898 586890 75454
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68058 -8694 68614
rect -8138 68058 30986 68614
rect 31542 68058 66986 68614
rect 67542 68058 102986 68614
rect 103542 68058 138986 68614
rect 139542 68058 174986 68614
rect 175542 68058 210986 68614
rect 211542 68058 246986 68614
rect 247542 68058 282986 68614
rect 283542 68058 318986 68614
rect 319542 68058 354986 68614
rect 355542 68058 390986 68614
rect 391542 68058 426986 68614
rect 427542 68058 462986 68614
rect 463542 68058 498986 68614
rect 499542 68058 534986 68614
rect 535542 68058 570986 68614
rect 571542 68058 592062 68614
rect 592618 68058 592650 68614
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64338 -6774 64894
rect -6218 64338 27266 64894
rect 27822 64338 63266 64894
rect 63822 64338 99266 64894
rect 99822 64338 135266 64894
rect 135822 64338 171266 64894
rect 171822 64338 207266 64894
rect 207822 64338 243266 64894
rect 243822 64338 279266 64894
rect 279822 64338 315266 64894
rect 315822 64338 351266 64894
rect 351822 64338 387266 64894
rect 387822 64338 423266 64894
rect 423822 64338 459266 64894
rect 459822 64338 495266 64894
rect 495822 64338 531266 64894
rect 531822 64338 567266 64894
rect 567822 64338 590142 64894
rect 590698 64338 590730 64894
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60618 -4854 61174
rect -4298 60618 23546 61174
rect 24102 60618 59546 61174
rect 60102 60618 95546 61174
rect 96102 60618 131546 61174
rect 132102 60618 167546 61174
rect 168102 60618 203546 61174
rect 204102 60618 239546 61174
rect 240102 60618 275546 61174
rect 276102 60618 311546 61174
rect 312102 60618 347546 61174
rect 348102 60618 383546 61174
rect 384102 60618 419546 61174
rect 420102 60618 455546 61174
rect 456102 60618 491546 61174
rect 492102 60618 527546 61174
rect 528102 60618 563546 61174
rect 564102 60618 588222 61174
rect 588778 60618 588810 61174
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 56898 -2934 57454
rect -2378 56898 19826 57454
rect 20382 56898 55826 57454
rect 56382 56898 91826 57454
rect 92382 56898 127826 57454
rect 128382 56898 163826 57454
rect 164382 56898 199826 57454
rect 200382 56898 235826 57454
rect 236382 56898 271826 57454
rect 272382 56898 307826 57454
rect 308382 56898 343826 57454
rect 344382 56898 379826 57454
rect 380382 56898 415826 57454
rect 416382 56898 451826 57454
rect 452382 56898 487826 57454
rect 488382 56898 523826 57454
rect 524382 56898 559826 57454
rect 560382 56898 586302 57454
rect 586858 56898 586890 57454
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50058 -7734 50614
rect -7178 50058 12986 50614
rect 13542 50058 48986 50614
rect 49542 50058 84986 50614
rect 85542 50058 120986 50614
rect 121542 50058 156986 50614
rect 157542 50058 192986 50614
rect 193542 50058 228986 50614
rect 229542 50058 264986 50614
rect 265542 50058 300986 50614
rect 301542 50058 336986 50614
rect 337542 50058 372986 50614
rect 373542 50058 408986 50614
rect 409542 50058 444986 50614
rect 445542 50058 480986 50614
rect 481542 50058 516986 50614
rect 517542 50058 552986 50614
rect 553542 50058 591102 50614
rect 591658 50058 592650 50614
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46338 -5814 46894
rect -5258 46338 9266 46894
rect 9822 46338 45266 46894
rect 45822 46338 81266 46894
rect 81822 46338 117266 46894
rect 117822 46338 153266 46894
rect 153822 46338 189266 46894
rect 189822 46338 225266 46894
rect 225822 46338 261266 46894
rect 261822 46338 297266 46894
rect 297822 46338 333266 46894
rect 333822 46338 369266 46894
rect 369822 46338 405266 46894
rect 405822 46338 441266 46894
rect 441822 46338 477266 46894
rect 477822 46338 513266 46894
rect 513822 46338 549266 46894
rect 549822 46338 589182 46894
rect 589738 46338 590730 46894
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42618 -3894 43174
rect -3338 42618 5546 43174
rect 6102 42618 41546 43174
rect 42102 42618 77546 43174
rect 78102 42618 113546 43174
rect 114102 42618 149546 43174
rect 150102 42618 185546 43174
rect 186102 42618 221546 43174
rect 222102 42618 257546 43174
rect 258102 42618 293546 43174
rect 294102 42618 329546 43174
rect 330102 42618 365546 43174
rect 366102 42618 401546 43174
rect 402102 42618 437546 43174
rect 438102 42618 473546 43174
rect 474102 42618 509546 43174
rect 510102 42618 545546 43174
rect 546102 42618 581546 43174
rect 582102 42618 587262 43174
rect 587818 42618 588810 43174
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 38898 -1974 39454
rect -1418 38898 1826 39454
rect 2382 38898 37826 39454
rect 38382 38898 73826 39454
rect 74382 38898 109826 39454
rect 110382 38898 145826 39454
rect 146382 38898 181826 39454
rect 182382 38898 217826 39454
rect 218382 38898 253826 39454
rect 254382 38898 289826 39454
rect 290382 38898 325826 39454
rect 326382 38898 361826 39454
rect 362382 38898 397826 39454
rect 398382 38898 433826 39454
rect 434382 38898 469826 39454
rect 470382 38898 505826 39454
rect 506382 38898 541826 39454
rect 542382 38898 577826 39454
rect 578382 38898 585342 39454
rect 585898 38898 586890 39454
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32058 -8694 32614
rect -8138 32058 30986 32614
rect 31542 32058 66986 32614
rect 67542 32058 102986 32614
rect 103542 32058 138986 32614
rect 139542 32058 174986 32614
rect 175542 32058 210986 32614
rect 211542 32058 246986 32614
rect 247542 32058 282986 32614
rect 283542 32058 318986 32614
rect 319542 32058 354986 32614
rect 355542 32058 390986 32614
rect 391542 32058 426986 32614
rect 427542 32058 462986 32614
rect 463542 32058 498986 32614
rect 499542 32058 534986 32614
rect 535542 32058 570986 32614
rect 571542 32058 592062 32614
rect 592618 32058 592650 32614
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28338 -6774 28894
rect -6218 28338 27266 28894
rect 27822 28338 63266 28894
rect 63822 28338 99266 28894
rect 99822 28338 135266 28894
rect 135822 28338 171266 28894
rect 171822 28338 207266 28894
rect 207822 28338 243266 28894
rect 243822 28338 279266 28894
rect 279822 28338 315266 28894
rect 315822 28338 351266 28894
rect 351822 28338 387266 28894
rect 387822 28338 423266 28894
rect 423822 28338 459266 28894
rect 459822 28338 495266 28894
rect 495822 28338 531266 28894
rect 531822 28338 567266 28894
rect 567822 28338 590142 28894
rect 590698 28338 590730 28894
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24618 -4854 25174
rect -4298 24618 23546 25174
rect 24102 24618 59546 25174
rect 60102 24618 95546 25174
rect 96102 24618 131546 25174
rect 132102 24618 167546 25174
rect 168102 24618 203546 25174
rect 204102 24618 239546 25174
rect 240102 24618 275546 25174
rect 276102 24618 311546 25174
rect 312102 24618 347546 25174
rect 348102 24618 383546 25174
rect 384102 24618 419546 25174
rect 420102 24618 455546 25174
rect 456102 24618 491546 25174
rect 492102 24618 527546 25174
rect 528102 24618 563546 25174
rect 564102 24618 588222 25174
rect 588778 24618 588810 25174
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 20898 -2934 21454
rect -2378 20898 19826 21454
rect 20382 20898 55826 21454
rect 56382 20898 91826 21454
rect 92382 20898 127826 21454
rect 128382 20898 163826 21454
rect 164382 20898 199826 21454
rect 200382 20898 235826 21454
rect 236382 20898 271826 21454
rect 272382 20898 307826 21454
rect 308382 20898 343826 21454
rect 344382 20898 379826 21454
rect 380382 20898 415826 21454
rect 416382 20898 451826 21454
rect 452382 20898 487826 21454
rect 488382 20898 523826 21454
rect 524382 20898 559826 21454
rect 560382 20898 586302 21454
rect 586858 20898 586890 21454
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14058 -7734 14614
rect -7178 14058 12986 14614
rect 13542 14058 48986 14614
rect 49542 14058 84986 14614
rect 85542 14058 120986 14614
rect 121542 14058 156986 14614
rect 157542 14058 192986 14614
rect 193542 14058 228986 14614
rect 229542 14058 264986 14614
rect 265542 14058 300986 14614
rect 301542 14058 336986 14614
rect 337542 14058 372986 14614
rect 373542 14058 408986 14614
rect 409542 14058 444986 14614
rect 445542 14058 480986 14614
rect 481542 14058 516986 14614
rect 517542 14058 552986 14614
rect 553542 14058 591102 14614
rect 591658 14058 592650 14614
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10338 -5814 10894
rect -5258 10338 9266 10894
rect 9822 10338 45266 10894
rect 45822 10338 81266 10894
rect 81822 10338 117266 10894
rect 117822 10338 153266 10894
rect 153822 10338 189266 10894
rect 189822 10338 225266 10894
rect 225822 10338 261266 10894
rect 261822 10338 297266 10894
rect 297822 10338 333266 10894
rect 333822 10338 369266 10894
rect 369822 10338 405266 10894
rect 405822 10338 441266 10894
rect 441822 10338 477266 10894
rect 477822 10338 513266 10894
rect 513822 10338 549266 10894
rect 549822 10338 589182 10894
rect 589738 10338 590730 10894
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6618 -3894 7174
rect -3338 6618 5546 7174
rect 6102 6618 41546 7174
rect 42102 6618 77546 7174
rect 78102 6618 113546 7174
rect 114102 6618 149546 7174
rect 150102 6618 185546 7174
rect 186102 6618 221546 7174
rect 222102 6618 257546 7174
rect 258102 6618 293546 7174
rect 294102 6618 329546 7174
rect 330102 6618 365546 7174
rect 366102 6618 401546 7174
rect 402102 6618 437546 7174
rect 438102 6618 473546 7174
rect 474102 6618 509546 7174
rect 510102 6618 545546 7174
rect 546102 6618 581546 7174
rect 582102 6618 587262 7174
rect 587818 6618 588810 7174
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 2898 -1974 3454
rect -1418 2898 1826 3454
rect 2382 2898 37826 3454
rect 38382 2898 73826 3454
rect 74382 2898 109826 3454
rect 110382 2898 145826 3454
rect 146382 2898 181826 3454
rect 182382 2898 217826 3454
rect 218382 2898 253826 3454
rect 254382 2898 289826 3454
rect 290382 2898 325826 3454
rect 326382 2898 361826 3454
rect 362382 2898 397826 3454
rect 398382 2898 433826 3454
rect 434382 2898 469826 3454
rect 470382 2898 505826 3454
rect 506382 2898 541826 3454
rect 542382 2898 577826 3454
rect 578382 2898 585342 3454
rect 585898 2898 586890 3454
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1826 -346
rect 2382 -902 37826 -346
rect 38382 -902 73826 -346
rect 74382 -902 109826 -346
rect 110382 -902 145826 -346
rect 146382 -902 181826 -346
rect 182382 -902 217826 -346
rect 218382 -902 253826 -346
rect 254382 -902 289826 -346
rect 290382 -902 325826 -346
rect 326382 -902 361826 -346
rect 362382 -902 397826 -346
rect 398382 -902 433826 -346
rect 434382 -902 469826 -346
rect 470382 -902 505826 -346
rect 506382 -902 541826 -346
rect 542382 -902 577826 -346
rect 578382 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 19826 -1306
rect 20382 -1862 55826 -1306
rect 56382 -1862 91826 -1306
rect 92382 -1862 127826 -1306
rect 128382 -1862 163826 -1306
rect 164382 -1862 199826 -1306
rect 200382 -1862 235826 -1306
rect 236382 -1862 271826 -1306
rect 272382 -1862 307826 -1306
rect 308382 -1862 343826 -1306
rect 344382 -1862 379826 -1306
rect 380382 -1862 415826 -1306
rect 416382 -1862 451826 -1306
rect 452382 -1862 487826 -1306
rect 488382 -1862 523826 -1306
rect 524382 -1862 559826 -1306
rect 560382 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 5546 -2266
rect 6102 -2822 41546 -2266
rect 42102 -2822 77546 -2266
rect 78102 -2822 113546 -2266
rect 114102 -2822 149546 -2266
rect 150102 -2822 185546 -2266
rect 186102 -2822 221546 -2266
rect 222102 -2822 257546 -2266
rect 258102 -2822 293546 -2266
rect 294102 -2822 329546 -2266
rect 330102 -2822 365546 -2266
rect 366102 -2822 401546 -2266
rect 402102 -2822 437546 -2266
rect 438102 -2822 473546 -2266
rect 474102 -2822 509546 -2266
rect 510102 -2822 545546 -2266
rect 546102 -2822 581546 -2266
rect 582102 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 23546 -3226
rect 24102 -3782 59546 -3226
rect 60102 -3782 95546 -3226
rect 96102 -3782 131546 -3226
rect 132102 -3782 167546 -3226
rect 168102 -3782 203546 -3226
rect 204102 -3782 239546 -3226
rect 240102 -3782 275546 -3226
rect 276102 -3782 311546 -3226
rect 312102 -3782 347546 -3226
rect 348102 -3782 383546 -3226
rect 384102 -3782 419546 -3226
rect 420102 -3782 455546 -3226
rect 456102 -3782 491546 -3226
rect 492102 -3782 527546 -3226
rect 528102 -3782 563546 -3226
rect 564102 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 9266 -4186
rect 9822 -4742 45266 -4186
rect 45822 -4742 81266 -4186
rect 81822 -4742 117266 -4186
rect 117822 -4742 153266 -4186
rect 153822 -4742 189266 -4186
rect 189822 -4742 225266 -4186
rect 225822 -4742 261266 -4186
rect 261822 -4742 297266 -4186
rect 297822 -4742 333266 -4186
rect 333822 -4742 369266 -4186
rect 369822 -4742 405266 -4186
rect 405822 -4742 441266 -4186
rect 441822 -4742 477266 -4186
rect 477822 -4742 513266 -4186
rect 513822 -4742 549266 -4186
rect 549822 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 27266 -5146
rect 27822 -5702 63266 -5146
rect 63822 -5702 99266 -5146
rect 99822 -5702 135266 -5146
rect 135822 -5702 171266 -5146
rect 171822 -5702 207266 -5146
rect 207822 -5702 243266 -5146
rect 243822 -5702 279266 -5146
rect 279822 -5702 315266 -5146
rect 315822 -5702 351266 -5146
rect 351822 -5702 387266 -5146
rect 387822 -5702 423266 -5146
rect 423822 -5702 459266 -5146
rect 459822 -5702 495266 -5146
rect 495822 -5702 531266 -5146
rect 531822 -5702 567266 -5146
rect 567822 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 12986 -6106
rect 13542 -6662 48986 -6106
rect 49542 -6662 84986 -6106
rect 85542 -6662 120986 -6106
rect 121542 -6662 156986 -6106
rect 157542 -6662 192986 -6106
rect 193542 -6662 228986 -6106
rect 229542 -6662 264986 -6106
rect 265542 -6662 300986 -6106
rect 301542 -6662 336986 -6106
rect 337542 -6662 372986 -6106
rect 373542 -6662 408986 -6106
rect 409542 -6662 444986 -6106
rect 445542 -6662 480986 -6106
rect 481542 -6662 516986 -6106
rect 517542 -6662 552986 -6106
rect 553542 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 30986 -7066
rect 31542 -7622 66986 -7066
rect 67542 -7622 102986 -7066
rect 103542 -7622 138986 -7066
rect 139542 -7622 174986 -7066
rect 175542 -7622 210986 -7066
rect 211542 -7622 246986 -7066
rect 247542 -7622 282986 -7066
rect 283542 -7622 318986 -7066
rect 319542 -7622 354986 -7066
rect 355542 -7622 390986 -7066
rect 391542 -7622 426986 -7066
rect 427542 -7622 462986 -7066
rect 463542 -7622 498986 -7066
rect 499542 -7622 534986 -7066
rect 535542 -7622 570986 -7066
rect 571542 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 235000 0 1 338000
box 198 0 199810 160000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 4 analog_io[0]
port 1 nsew
rlabel metal2 s 446098 703520 446210 704960 4 analog_io[10]
port 2 nsew
rlabel metal2 s 381146 703520 381258 704960 4 analog_io[11]
port 3 nsew
rlabel metal2 s 316286 703520 316398 704960 4 analog_io[12]
port 4 nsew
rlabel metal2 s 251426 703520 251538 704960 4 analog_io[13]
port 5 nsew
rlabel metal2 s 186474 703520 186586 704960 4 analog_io[14]
port 6 nsew
rlabel metal2 s 121614 703520 121726 704960 4 analog_io[15]
port 7 nsew
rlabel metal2 s 56754 703520 56866 704960 4 analog_io[16]
port 8 nsew
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew
rlabel metal3 s 583520 338452 584960 338692 4 analog_io[1]
port 12 nsew
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew
rlabel metal3 s 583520 391628 584960 391868 4 analog_io[2]
port 22 nsew
rlabel metal3 s 583520 444668 584960 444908 4 analog_io[3]
port 23 nsew
rlabel metal3 s 583520 497844 584960 498084 4 analog_io[4]
port 24 nsew
rlabel metal3 s 583520 551020 584960 551260 4 analog_io[5]
port 25 nsew
rlabel metal3 s 583520 604060 584960 604300 4 analog_io[6]
port 26 nsew
rlabel metal3 s 583520 657236 584960 657476 4 analog_io[7]
port 27 nsew
rlabel metal2 s 575818 703520 575930 704960 4 analog_io[8]
port 28 nsew
rlabel metal2 s 510958 703520 511070 704960 4 analog_io[9]
port 29 nsew
rlabel metal3 s 583520 6476 584960 6716 4 io_in[0]
port 30 nsew
rlabel metal3 s 583520 457996 584960 458236 4 io_in[10]
port 31 nsew
rlabel metal3 s 583520 511172 584960 511412 4 io_in[11]
port 32 nsew
rlabel metal3 s 583520 564212 584960 564452 4 io_in[12]
port 33 nsew
rlabel metal3 s 583520 617388 584960 617628 4 io_in[13]
port 34 nsew
rlabel metal3 s 583520 670564 584960 670804 4 io_in[14]
port 35 nsew
rlabel metal2 s 559626 703520 559738 704960 4 io_in[15]
port 36 nsew
rlabel metal2 s 494766 703520 494878 704960 4 io_in[16]
port 37 nsew
rlabel metal2 s 429814 703520 429926 704960 4 io_in[17]
port 38 nsew
rlabel metal2 s 364954 703520 365066 704960 4 io_in[18]
port 39 nsew
rlabel metal2 s 300094 703520 300206 704960 4 io_in[19]
port 40 nsew
rlabel metal3 s 583520 46188 584960 46428 4 io_in[1]
port 41 nsew
rlabel metal2 s 235142 703520 235254 704960 4 io_in[20]
port 42 nsew
rlabel metal2 s 170282 703520 170394 704960 4 io_in[21]
port 43 nsew
rlabel metal2 s 105422 703520 105534 704960 4 io_in[22]
port 44 nsew
rlabel metal2 s 40470 703520 40582 704960 4 io_in[23]
port 45 nsew
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew
rlabel metal3 s 583520 86036 584960 86276 4 io_in[2]
port 52 nsew
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew
rlabel metal3 s 583520 125884 584960 126124 4 io_in[3]
port 61 nsew
rlabel metal3 s 583520 165732 584960 165972 4 io_in[4]
port 62 nsew
rlabel metal3 s 583520 205580 584960 205820 4 io_in[5]
port 63 nsew
rlabel metal3 s 583520 245428 584960 245668 4 io_in[6]
port 64 nsew
rlabel metal3 s 583520 298604 584960 298844 4 io_in[7]
port 65 nsew
rlabel metal3 s 583520 351780 584960 352020 4 io_in[8]
port 66 nsew
rlabel metal3 s 583520 404820 584960 405060 4 io_in[9]
port 67 nsew
rlabel metal3 s 583520 32996 584960 33236 4 io_oeb[0]
port 68 nsew
rlabel metal3 s 583520 484516 584960 484756 4 io_oeb[10]
port 69 nsew
rlabel metal3 s 583520 537692 584960 537932 4 io_oeb[11]
port 70 nsew
rlabel metal3 s 583520 590868 584960 591108 4 io_oeb[12]
port 71 nsew
rlabel metal3 s 583520 643908 584960 644148 4 io_oeb[13]
port 72 nsew
rlabel metal3 s 583520 697084 584960 697324 4 io_oeb[14]
port 73 nsew
rlabel metal2 s 527150 703520 527262 704960 4 io_oeb[15]
port 74 nsew
rlabel metal2 s 462290 703520 462402 704960 4 io_oeb[16]
port 75 nsew
rlabel metal2 s 397430 703520 397542 704960 4 io_oeb[17]
port 76 nsew
rlabel metal2 s 332478 703520 332590 704960 4 io_oeb[18]
port 77 nsew
rlabel metal2 s 267618 703520 267730 704960 4 io_oeb[19]
port 78 nsew
rlabel metal3 s 583520 72844 584960 73084 4 io_oeb[1]
port 79 nsew
rlabel metal2 s 202758 703520 202870 704960 4 io_oeb[20]
port 80 nsew
rlabel metal2 s 137806 703520 137918 704960 4 io_oeb[21]
port 81 nsew
rlabel metal2 s 72946 703520 73058 704960 4 io_oeb[22]
port 82 nsew
rlabel metal2 s 8086 703520 8198 704960 4 io_oeb[23]
port 83 nsew
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew
rlabel metal3 s 583520 112692 584960 112932 4 io_oeb[2]
port 90 nsew
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew
rlabel metal3 s 583520 152540 584960 152780 4 io_oeb[3]
port 99 nsew
rlabel metal3 s 583520 192388 584960 192628 4 io_oeb[4]
port 100 nsew
rlabel metal3 s 583520 232236 584960 232476 4 io_oeb[5]
port 101 nsew
rlabel metal3 s 583520 272084 584960 272324 4 io_oeb[6]
port 102 nsew
rlabel metal3 s 583520 325124 584960 325364 4 io_oeb[7]
port 103 nsew
rlabel metal3 s 583520 378300 584960 378540 4 io_oeb[8]
port 104 nsew
rlabel metal3 s 583520 431476 584960 431716 4 io_oeb[9]
port 105 nsew
rlabel metal3 s 583520 19668 584960 19908 4 io_out[0]
port 106 nsew
rlabel metal3 s 583520 471324 584960 471564 4 io_out[10]
port 107 nsew
rlabel metal3 s 583520 524364 584960 524604 4 io_out[11]
port 108 nsew
rlabel metal3 s 583520 577540 584960 577780 4 io_out[12]
port 109 nsew
rlabel metal3 s 583520 630716 584960 630956 4 io_out[13]
port 110 nsew
rlabel metal3 s 583520 683756 584960 683996 4 io_out[14]
port 111 nsew
rlabel metal2 s 543434 703520 543546 704960 4 io_out[15]
port 112 nsew
rlabel metal2 s 478482 703520 478594 704960 4 io_out[16]
port 113 nsew
rlabel metal2 s 413622 703520 413734 704960 4 io_out[17]
port 114 nsew
rlabel metal2 s 348762 703520 348874 704960 4 io_out[18]
port 115 nsew
rlabel metal2 s 283810 703520 283922 704960 4 io_out[19]
port 116 nsew
rlabel metal3 s 583520 59516 584960 59756 4 io_out[1]
port 117 nsew
rlabel metal2 s 218950 703520 219062 704960 4 io_out[20]
port 118 nsew
rlabel metal2 s 154090 703520 154202 704960 4 io_out[21]
port 119 nsew
rlabel metal2 s 89138 703520 89250 704960 4 io_out[22]
port 120 nsew
rlabel metal2 s 24278 703520 24390 704960 4 io_out[23]
port 121 nsew
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew
rlabel metal3 s 583520 99364 584960 99604 4 io_out[2]
port 128 nsew
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew
rlabel metal3 s 583520 139212 584960 139452 4 io_out[3]
port 137 nsew
rlabel metal3 s 583520 179060 584960 179300 4 io_out[4]
port 138 nsew
rlabel metal3 s 583520 218908 584960 219148 4 io_out[5]
port 139 nsew
rlabel metal3 s 583520 258756 584960 258996 4 io_out[6]
port 140 nsew
rlabel metal3 s 583520 311932 584960 312172 4 io_out[7]
port 141 nsew
rlabel metal3 s 583520 364972 584960 365212 4 io_out[8]
port 142 nsew
rlabel metal3 s 583520 418148 584960 418388 4 io_out[9]
port 143 nsew
rlabel metal2 s 125846 -960 125958 480 4 la_data_in[0]
port 144 nsew
rlabel metal2 s 480506 -960 480618 480 4 la_data_in[100]
port 145 nsew
rlabel metal2 s 484002 -960 484114 480 4 la_data_in[101]
port 146 nsew
rlabel metal2 s 487590 -960 487702 480 4 la_data_in[102]
port 147 nsew
rlabel metal2 s 491086 -960 491198 480 4 la_data_in[103]
port 148 nsew
rlabel metal2 s 494674 -960 494786 480 4 la_data_in[104]
port 149 nsew
rlabel metal2 s 498170 -960 498282 480 4 la_data_in[105]
port 150 nsew
rlabel metal2 s 501758 -960 501870 480 4 la_data_in[106]
port 151 nsew
rlabel metal2 s 505346 -960 505458 480 4 la_data_in[107]
port 152 nsew
rlabel metal2 s 508842 -960 508954 480 4 la_data_in[108]
port 153 nsew
rlabel metal2 s 512430 -960 512542 480 4 la_data_in[109]
port 154 nsew
rlabel metal2 s 161266 -960 161378 480 4 la_data_in[10]
port 155 nsew
rlabel metal2 s 515926 -960 516038 480 4 la_data_in[110]
port 156 nsew
rlabel metal2 s 519514 -960 519626 480 4 la_data_in[111]
port 157 nsew
rlabel metal2 s 523010 -960 523122 480 4 la_data_in[112]
port 158 nsew
rlabel metal2 s 526598 -960 526710 480 4 la_data_in[113]
port 159 nsew
rlabel metal2 s 530094 -960 530206 480 4 la_data_in[114]
port 160 nsew
rlabel metal2 s 533682 -960 533794 480 4 la_data_in[115]
port 161 nsew
rlabel metal2 s 537178 -960 537290 480 4 la_data_in[116]
port 162 nsew
rlabel metal2 s 540766 -960 540878 480 4 la_data_in[117]
port 163 nsew
rlabel metal2 s 544354 -960 544466 480 4 la_data_in[118]
port 164 nsew
rlabel metal2 s 547850 -960 547962 480 4 la_data_in[119]
port 165 nsew
rlabel metal2 s 164854 -960 164966 480 4 la_data_in[11]
port 166 nsew
rlabel metal2 s 551438 -960 551550 480 4 la_data_in[120]
port 167 nsew
rlabel metal2 s 554934 -960 555046 480 4 la_data_in[121]
port 168 nsew
rlabel metal2 s 558522 -960 558634 480 4 la_data_in[122]
port 169 nsew
rlabel metal2 s 562018 -960 562130 480 4 la_data_in[123]
port 170 nsew
rlabel metal2 s 565606 -960 565718 480 4 la_data_in[124]
port 171 nsew
rlabel metal2 s 569102 -960 569214 480 4 la_data_in[125]
port 172 nsew
rlabel metal2 s 572690 -960 572802 480 4 la_data_in[126]
port 173 nsew
rlabel metal2 s 576278 -960 576390 480 4 la_data_in[127]
port 174 nsew
rlabel metal2 s 168350 -960 168462 480 4 la_data_in[12]
port 175 nsew
rlabel metal2 s 171938 -960 172050 480 4 la_data_in[13]
port 176 nsew
rlabel metal2 s 175434 -960 175546 480 4 la_data_in[14]
port 177 nsew
rlabel metal2 s 179022 -960 179134 480 4 la_data_in[15]
port 178 nsew
rlabel metal2 s 182518 -960 182630 480 4 la_data_in[16]
port 179 nsew
rlabel metal2 s 186106 -960 186218 480 4 la_data_in[17]
port 180 nsew
rlabel metal2 s 189694 -960 189806 480 4 la_data_in[18]
port 181 nsew
rlabel metal2 s 193190 -960 193302 480 4 la_data_in[19]
port 182 nsew
rlabel metal2 s 129342 -960 129454 480 4 la_data_in[1]
port 183 nsew
rlabel metal2 s 196778 -960 196890 480 4 la_data_in[20]
port 184 nsew
rlabel metal2 s 200274 -960 200386 480 4 la_data_in[21]
port 185 nsew
rlabel metal2 s 203862 -960 203974 480 4 la_data_in[22]
port 186 nsew
rlabel metal2 s 207358 -960 207470 480 4 la_data_in[23]
port 187 nsew
rlabel metal2 s 210946 -960 211058 480 4 la_data_in[24]
port 188 nsew
rlabel metal2 s 214442 -960 214554 480 4 la_data_in[25]
port 189 nsew
rlabel metal2 s 218030 -960 218142 480 4 la_data_in[26]
port 190 nsew
rlabel metal2 s 221526 -960 221638 480 4 la_data_in[27]
port 191 nsew
rlabel metal2 s 225114 -960 225226 480 4 la_data_in[28]
port 192 nsew
rlabel metal2 s 228702 -960 228814 480 4 la_data_in[29]
port 193 nsew
rlabel metal2 s 132930 -960 133042 480 4 la_data_in[2]
port 194 nsew
rlabel metal2 s 232198 -960 232310 480 4 la_data_in[30]
port 195 nsew
rlabel metal2 s 235786 -960 235898 480 4 la_data_in[31]
port 196 nsew
rlabel metal2 s 239282 -960 239394 480 4 la_data_in[32]
port 197 nsew
rlabel metal2 s 242870 -960 242982 480 4 la_data_in[33]
port 198 nsew
rlabel metal2 s 246366 -960 246478 480 4 la_data_in[34]
port 199 nsew
rlabel metal2 s 249954 -960 250066 480 4 la_data_in[35]
port 200 nsew
rlabel metal2 s 253450 -960 253562 480 4 la_data_in[36]
port 201 nsew
rlabel metal2 s 257038 -960 257150 480 4 la_data_in[37]
port 202 nsew
rlabel metal2 s 260626 -960 260738 480 4 la_data_in[38]
port 203 nsew
rlabel metal2 s 264122 -960 264234 480 4 la_data_in[39]
port 204 nsew
rlabel metal2 s 136426 -960 136538 480 4 la_data_in[3]
port 205 nsew
rlabel metal2 s 267710 -960 267822 480 4 la_data_in[40]
port 206 nsew
rlabel metal2 s 271206 -960 271318 480 4 la_data_in[41]
port 207 nsew
rlabel metal2 s 274794 -960 274906 480 4 la_data_in[42]
port 208 nsew
rlabel metal2 s 278290 -960 278402 480 4 la_data_in[43]
port 209 nsew
rlabel metal2 s 281878 -960 281990 480 4 la_data_in[44]
port 210 nsew
rlabel metal2 s 285374 -960 285486 480 4 la_data_in[45]
port 211 nsew
rlabel metal2 s 288962 -960 289074 480 4 la_data_in[46]
port 212 nsew
rlabel metal2 s 292550 -960 292662 480 4 la_data_in[47]
port 213 nsew
rlabel metal2 s 296046 -960 296158 480 4 la_data_in[48]
port 214 nsew
rlabel metal2 s 299634 -960 299746 480 4 la_data_in[49]
port 215 nsew
rlabel metal2 s 140014 -960 140126 480 4 la_data_in[4]
port 216 nsew
rlabel metal2 s 303130 -960 303242 480 4 la_data_in[50]
port 217 nsew
rlabel metal2 s 306718 -960 306830 480 4 la_data_in[51]
port 218 nsew
rlabel metal2 s 310214 -960 310326 480 4 la_data_in[52]
port 219 nsew
rlabel metal2 s 313802 -960 313914 480 4 la_data_in[53]
port 220 nsew
rlabel metal2 s 317298 -960 317410 480 4 la_data_in[54]
port 221 nsew
rlabel metal2 s 320886 -960 320998 480 4 la_data_in[55]
port 222 nsew
rlabel metal2 s 324382 -960 324494 480 4 la_data_in[56]
port 223 nsew
rlabel metal2 s 327970 -960 328082 480 4 la_data_in[57]
port 224 nsew
rlabel metal2 s 331558 -960 331670 480 4 la_data_in[58]
port 225 nsew
rlabel metal2 s 335054 -960 335166 480 4 la_data_in[59]
port 226 nsew
rlabel metal2 s 143510 -960 143622 480 4 la_data_in[5]
port 227 nsew
rlabel metal2 s 338642 -960 338754 480 4 la_data_in[60]
port 228 nsew
rlabel metal2 s 342138 -960 342250 480 4 la_data_in[61]
port 229 nsew
rlabel metal2 s 345726 -960 345838 480 4 la_data_in[62]
port 230 nsew
rlabel metal2 s 349222 -960 349334 480 4 la_data_in[63]
port 231 nsew
rlabel metal2 s 352810 -960 352922 480 4 la_data_in[64]
port 232 nsew
rlabel metal2 s 356306 -960 356418 480 4 la_data_in[65]
port 233 nsew
rlabel metal2 s 359894 -960 360006 480 4 la_data_in[66]
port 234 nsew
rlabel metal2 s 363482 -960 363594 480 4 la_data_in[67]
port 235 nsew
rlabel metal2 s 366978 -960 367090 480 4 la_data_in[68]
port 236 nsew
rlabel metal2 s 370566 -960 370678 480 4 la_data_in[69]
port 237 nsew
rlabel metal2 s 147098 -960 147210 480 4 la_data_in[6]
port 238 nsew
rlabel metal2 s 374062 -960 374174 480 4 la_data_in[70]
port 239 nsew
rlabel metal2 s 377650 -960 377762 480 4 la_data_in[71]
port 240 nsew
rlabel metal2 s 381146 -960 381258 480 4 la_data_in[72]
port 241 nsew
rlabel metal2 s 384734 -960 384846 480 4 la_data_in[73]
port 242 nsew
rlabel metal2 s 388230 -960 388342 480 4 la_data_in[74]
port 243 nsew
rlabel metal2 s 391818 -960 391930 480 4 la_data_in[75]
port 244 nsew
rlabel metal2 s 395314 -960 395426 480 4 la_data_in[76]
port 245 nsew
rlabel metal2 s 398902 -960 399014 480 4 la_data_in[77]
port 246 nsew
rlabel metal2 s 402490 -960 402602 480 4 la_data_in[78]
port 247 nsew
rlabel metal2 s 405986 -960 406098 480 4 la_data_in[79]
port 248 nsew
rlabel metal2 s 150594 -960 150706 480 4 la_data_in[7]
port 249 nsew
rlabel metal2 s 409574 -960 409686 480 4 la_data_in[80]
port 250 nsew
rlabel metal2 s 413070 -960 413182 480 4 la_data_in[81]
port 251 nsew
rlabel metal2 s 416658 -960 416770 480 4 la_data_in[82]
port 252 nsew
rlabel metal2 s 420154 -960 420266 480 4 la_data_in[83]
port 253 nsew
rlabel metal2 s 423742 -960 423854 480 4 la_data_in[84]
port 254 nsew
rlabel metal2 s 427238 -960 427350 480 4 la_data_in[85]
port 255 nsew
rlabel metal2 s 430826 -960 430938 480 4 la_data_in[86]
port 256 nsew
rlabel metal2 s 434414 -960 434526 480 4 la_data_in[87]
port 257 nsew
rlabel metal2 s 437910 -960 438022 480 4 la_data_in[88]
port 258 nsew
rlabel metal2 s 441498 -960 441610 480 4 la_data_in[89]
port 259 nsew
rlabel metal2 s 154182 -960 154294 480 4 la_data_in[8]
port 260 nsew
rlabel metal2 s 444994 -960 445106 480 4 la_data_in[90]
port 261 nsew
rlabel metal2 s 448582 -960 448694 480 4 la_data_in[91]
port 262 nsew
rlabel metal2 s 452078 -960 452190 480 4 la_data_in[92]
port 263 nsew
rlabel metal2 s 455666 -960 455778 480 4 la_data_in[93]
port 264 nsew
rlabel metal2 s 459162 -960 459274 480 4 la_data_in[94]
port 265 nsew
rlabel metal2 s 462750 -960 462862 480 4 la_data_in[95]
port 266 nsew
rlabel metal2 s 466246 -960 466358 480 4 la_data_in[96]
port 267 nsew
rlabel metal2 s 469834 -960 469946 480 4 la_data_in[97]
port 268 nsew
rlabel metal2 s 473422 -960 473534 480 4 la_data_in[98]
port 269 nsew
rlabel metal2 s 476918 -960 477030 480 4 la_data_in[99]
port 270 nsew
rlabel metal2 s 157770 -960 157882 480 4 la_data_in[9]
port 271 nsew
rlabel metal2 s 126950 -960 127062 480 4 la_data_out[0]
port 272 nsew
rlabel metal2 s 481702 -960 481814 480 4 la_data_out[100]
port 273 nsew
rlabel metal2 s 485198 -960 485310 480 4 la_data_out[101]
port 274 nsew
rlabel metal2 s 488786 -960 488898 480 4 la_data_out[102]
port 275 nsew
rlabel metal2 s 492282 -960 492394 480 4 la_data_out[103]
port 276 nsew
rlabel metal2 s 495870 -960 495982 480 4 la_data_out[104]
port 277 nsew
rlabel metal2 s 499366 -960 499478 480 4 la_data_out[105]
port 278 nsew
rlabel metal2 s 502954 -960 503066 480 4 la_data_out[106]
port 279 nsew
rlabel metal2 s 506450 -960 506562 480 4 la_data_out[107]
port 280 nsew
rlabel metal2 s 510038 -960 510150 480 4 la_data_out[108]
port 281 nsew
rlabel metal2 s 513534 -960 513646 480 4 la_data_out[109]
port 282 nsew
rlabel metal2 s 162462 -960 162574 480 4 la_data_out[10]
port 283 nsew
rlabel metal2 s 517122 -960 517234 480 4 la_data_out[110]
port 284 nsew
rlabel metal2 s 520710 -960 520822 480 4 la_data_out[111]
port 285 nsew
rlabel metal2 s 524206 -960 524318 480 4 la_data_out[112]
port 286 nsew
rlabel metal2 s 527794 -960 527906 480 4 la_data_out[113]
port 287 nsew
rlabel metal2 s 531290 -960 531402 480 4 la_data_out[114]
port 288 nsew
rlabel metal2 s 534878 -960 534990 480 4 la_data_out[115]
port 289 nsew
rlabel metal2 s 538374 -960 538486 480 4 la_data_out[116]
port 290 nsew
rlabel metal2 s 541962 -960 542074 480 4 la_data_out[117]
port 291 nsew
rlabel metal2 s 545458 -960 545570 480 4 la_data_out[118]
port 292 nsew
rlabel metal2 s 549046 -960 549158 480 4 la_data_out[119]
port 293 nsew
rlabel metal2 s 166050 -960 166162 480 4 la_data_out[11]
port 294 nsew
rlabel metal2 s 552634 -960 552746 480 4 la_data_out[120]
port 295 nsew
rlabel metal2 s 556130 -960 556242 480 4 la_data_out[121]
port 296 nsew
rlabel metal2 s 559718 -960 559830 480 4 la_data_out[122]
port 297 nsew
rlabel metal2 s 563214 -960 563326 480 4 la_data_out[123]
port 298 nsew
rlabel metal2 s 566802 -960 566914 480 4 la_data_out[124]
port 299 nsew
rlabel metal2 s 570298 -960 570410 480 4 la_data_out[125]
port 300 nsew
rlabel metal2 s 573886 -960 573998 480 4 la_data_out[126]
port 301 nsew
rlabel metal2 s 577382 -960 577494 480 4 la_data_out[127]
port 302 nsew
rlabel metal2 s 169546 -960 169658 480 4 la_data_out[12]
port 303 nsew
rlabel metal2 s 173134 -960 173246 480 4 la_data_out[13]
port 304 nsew
rlabel metal2 s 176630 -960 176742 480 4 la_data_out[14]
port 305 nsew
rlabel metal2 s 180218 -960 180330 480 4 la_data_out[15]
port 306 nsew
rlabel metal2 s 183714 -960 183826 480 4 la_data_out[16]
port 307 nsew
rlabel metal2 s 187302 -960 187414 480 4 la_data_out[17]
port 308 nsew
rlabel metal2 s 190798 -960 190910 480 4 la_data_out[18]
port 309 nsew
rlabel metal2 s 194386 -960 194498 480 4 la_data_out[19]
port 310 nsew
rlabel metal2 s 130538 -960 130650 480 4 la_data_out[1]
port 311 nsew
rlabel metal2 s 197882 -960 197994 480 4 la_data_out[20]
port 312 nsew
rlabel metal2 s 201470 -960 201582 480 4 la_data_out[21]
port 313 nsew
rlabel metal2 s 205058 -960 205170 480 4 la_data_out[22]
port 314 nsew
rlabel metal2 s 208554 -960 208666 480 4 la_data_out[23]
port 315 nsew
rlabel metal2 s 212142 -960 212254 480 4 la_data_out[24]
port 316 nsew
rlabel metal2 s 215638 -960 215750 480 4 la_data_out[25]
port 317 nsew
rlabel metal2 s 219226 -960 219338 480 4 la_data_out[26]
port 318 nsew
rlabel metal2 s 222722 -960 222834 480 4 la_data_out[27]
port 319 nsew
rlabel metal2 s 226310 -960 226422 480 4 la_data_out[28]
port 320 nsew
rlabel metal2 s 229806 -960 229918 480 4 la_data_out[29]
port 321 nsew
rlabel metal2 s 134126 -960 134238 480 4 la_data_out[2]
port 322 nsew
rlabel metal2 s 233394 -960 233506 480 4 la_data_out[30]
port 323 nsew
rlabel metal2 s 236982 -960 237094 480 4 la_data_out[31]
port 324 nsew
rlabel metal2 s 240478 -960 240590 480 4 la_data_out[32]
port 325 nsew
rlabel metal2 s 244066 -960 244178 480 4 la_data_out[33]
port 326 nsew
rlabel metal2 s 247562 -960 247674 480 4 la_data_out[34]
port 327 nsew
rlabel metal2 s 251150 -960 251262 480 4 la_data_out[35]
port 328 nsew
rlabel metal2 s 254646 -960 254758 480 4 la_data_out[36]
port 329 nsew
rlabel metal2 s 258234 -960 258346 480 4 la_data_out[37]
port 330 nsew
rlabel metal2 s 261730 -960 261842 480 4 la_data_out[38]
port 331 nsew
rlabel metal2 s 265318 -960 265430 480 4 la_data_out[39]
port 332 nsew
rlabel metal2 s 137622 -960 137734 480 4 la_data_out[3]
port 333 nsew
rlabel metal2 s 268814 -960 268926 480 4 la_data_out[40]
port 334 nsew
rlabel metal2 s 272402 -960 272514 480 4 la_data_out[41]
port 335 nsew
rlabel metal2 s 275990 -960 276102 480 4 la_data_out[42]
port 336 nsew
rlabel metal2 s 279486 -960 279598 480 4 la_data_out[43]
port 337 nsew
rlabel metal2 s 283074 -960 283186 480 4 la_data_out[44]
port 338 nsew
rlabel metal2 s 286570 -960 286682 480 4 la_data_out[45]
port 339 nsew
rlabel metal2 s 290158 -960 290270 480 4 la_data_out[46]
port 340 nsew
rlabel metal2 s 293654 -960 293766 480 4 la_data_out[47]
port 341 nsew
rlabel metal2 s 297242 -960 297354 480 4 la_data_out[48]
port 342 nsew
rlabel metal2 s 300738 -960 300850 480 4 la_data_out[49]
port 343 nsew
rlabel metal2 s 141210 -960 141322 480 4 la_data_out[4]
port 344 nsew
rlabel metal2 s 304326 -960 304438 480 4 la_data_out[50]
port 345 nsew
rlabel metal2 s 307914 -960 308026 480 4 la_data_out[51]
port 346 nsew
rlabel metal2 s 311410 -960 311522 480 4 la_data_out[52]
port 347 nsew
rlabel metal2 s 314998 -960 315110 480 4 la_data_out[53]
port 348 nsew
rlabel metal2 s 318494 -960 318606 480 4 la_data_out[54]
port 349 nsew
rlabel metal2 s 322082 -960 322194 480 4 la_data_out[55]
port 350 nsew
rlabel metal2 s 325578 -960 325690 480 4 la_data_out[56]
port 351 nsew
rlabel metal2 s 329166 -960 329278 480 4 la_data_out[57]
port 352 nsew
rlabel metal2 s 332662 -960 332774 480 4 la_data_out[58]
port 353 nsew
rlabel metal2 s 336250 -960 336362 480 4 la_data_out[59]
port 354 nsew
rlabel metal2 s 144706 -960 144818 480 4 la_data_out[5]
port 355 nsew
rlabel metal2 s 339838 -960 339950 480 4 la_data_out[60]
port 356 nsew
rlabel metal2 s 343334 -960 343446 480 4 la_data_out[61]
port 357 nsew
rlabel metal2 s 346922 -960 347034 480 4 la_data_out[62]
port 358 nsew
rlabel metal2 s 350418 -960 350530 480 4 la_data_out[63]
port 359 nsew
rlabel metal2 s 354006 -960 354118 480 4 la_data_out[64]
port 360 nsew
rlabel metal2 s 357502 -960 357614 480 4 la_data_out[65]
port 361 nsew
rlabel metal2 s 361090 -960 361202 480 4 la_data_out[66]
port 362 nsew
rlabel metal2 s 364586 -960 364698 480 4 la_data_out[67]
port 363 nsew
rlabel metal2 s 368174 -960 368286 480 4 la_data_out[68]
port 364 nsew
rlabel metal2 s 371670 -960 371782 480 4 la_data_out[69]
port 365 nsew
rlabel metal2 s 148294 -960 148406 480 4 la_data_out[6]
port 366 nsew
rlabel metal2 s 375258 -960 375370 480 4 la_data_out[70]
port 367 nsew
rlabel metal2 s 378846 -960 378958 480 4 la_data_out[71]
port 368 nsew
rlabel metal2 s 382342 -960 382454 480 4 la_data_out[72]
port 369 nsew
rlabel metal2 s 385930 -960 386042 480 4 la_data_out[73]
port 370 nsew
rlabel metal2 s 389426 -960 389538 480 4 la_data_out[74]
port 371 nsew
rlabel metal2 s 393014 -960 393126 480 4 la_data_out[75]
port 372 nsew
rlabel metal2 s 396510 -960 396622 480 4 la_data_out[76]
port 373 nsew
rlabel metal2 s 400098 -960 400210 480 4 la_data_out[77]
port 374 nsew
rlabel metal2 s 403594 -960 403706 480 4 la_data_out[78]
port 375 nsew
rlabel metal2 s 407182 -960 407294 480 4 la_data_out[79]
port 376 nsew
rlabel metal2 s 151790 -960 151902 480 4 la_data_out[7]
port 377 nsew
rlabel metal2 s 410770 -960 410882 480 4 la_data_out[80]
port 378 nsew
rlabel metal2 s 414266 -960 414378 480 4 la_data_out[81]
port 379 nsew
rlabel metal2 s 417854 -960 417966 480 4 la_data_out[82]
port 380 nsew
rlabel metal2 s 421350 -960 421462 480 4 la_data_out[83]
port 381 nsew
rlabel metal2 s 424938 -960 425050 480 4 la_data_out[84]
port 382 nsew
rlabel metal2 s 428434 -960 428546 480 4 la_data_out[85]
port 383 nsew
rlabel metal2 s 432022 -960 432134 480 4 la_data_out[86]
port 384 nsew
rlabel metal2 s 435518 -960 435630 480 4 la_data_out[87]
port 385 nsew
rlabel metal2 s 439106 -960 439218 480 4 la_data_out[88]
port 386 nsew
rlabel metal2 s 442602 -960 442714 480 4 la_data_out[89]
port 387 nsew
rlabel metal2 s 155378 -960 155490 480 4 la_data_out[8]
port 388 nsew
rlabel metal2 s 446190 -960 446302 480 4 la_data_out[90]
port 389 nsew
rlabel metal2 s 449778 -960 449890 480 4 la_data_out[91]
port 390 nsew
rlabel metal2 s 453274 -960 453386 480 4 la_data_out[92]
port 391 nsew
rlabel metal2 s 456862 -960 456974 480 4 la_data_out[93]
port 392 nsew
rlabel metal2 s 460358 -960 460470 480 4 la_data_out[94]
port 393 nsew
rlabel metal2 s 463946 -960 464058 480 4 la_data_out[95]
port 394 nsew
rlabel metal2 s 467442 -960 467554 480 4 la_data_out[96]
port 395 nsew
rlabel metal2 s 471030 -960 471142 480 4 la_data_out[97]
port 396 nsew
rlabel metal2 s 474526 -960 474638 480 4 la_data_out[98]
port 397 nsew
rlabel metal2 s 478114 -960 478226 480 4 la_data_out[99]
port 398 nsew
rlabel metal2 s 158874 -960 158986 480 4 la_data_out[9]
port 399 nsew
rlabel metal2 s 128146 -960 128258 480 4 la_oenb[0]
port 400 nsew
rlabel metal2 s 482806 -960 482918 480 4 la_oenb[100]
port 401 nsew
rlabel metal2 s 486394 -960 486506 480 4 la_oenb[101]
port 402 nsew
rlabel metal2 s 489890 -960 490002 480 4 la_oenb[102]
port 403 nsew
rlabel metal2 s 493478 -960 493590 480 4 la_oenb[103]
port 404 nsew
rlabel metal2 s 497066 -960 497178 480 4 la_oenb[104]
port 405 nsew
rlabel metal2 s 500562 -960 500674 480 4 la_oenb[105]
port 406 nsew
rlabel metal2 s 504150 -960 504262 480 4 la_oenb[106]
port 407 nsew
rlabel metal2 s 507646 -960 507758 480 4 la_oenb[107]
port 408 nsew
rlabel metal2 s 511234 -960 511346 480 4 la_oenb[108]
port 409 nsew
rlabel metal2 s 514730 -960 514842 480 4 la_oenb[109]
port 410 nsew
rlabel metal2 s 163658 -960 163770 480 4 la_oenb[10]
port 411 nsew
rlabel metal2 s 518318 -960 518430 480 4 la_oenb[110]
port 412 nsew
rlabel metal2 s 521814 -960 521926 480 4 la_oenb[111]
port 413 nsew
rlabel metal2 s 525402 -960 525514 480 4 la_oenb[112]
port 414 nsew
rlabel metal2 s 528990 -960 529102 480 4 la_oenb[113]
port 415 nsew
rlabel metal2 s 532486 -960 532598 480 4 la_oenb[114]
port 416 nsew
rlabel metal2 s 536074 -960 536186 480 4 la_oenb[115]
port 417 nsew
rlabel metal2 s 539570 -960 539682 480 4 la_oenb[116]
port 418 nsew
rlabel metal2 s 543158 -960 543270 480 4 la_oenb[117]
port 419 nsew
rlabel metal2 s 546654 -960 546766 480 4 la_oenb[118]
port 420 nsew
rlabel metal2 s 550242 -960 550354 480 4 la_oenb[119]
port 421 nsew
rlabel metal2 s 167154 -960 167266 480 4 la_oenb[11]
port 422 nsew
rlabel metal2 s 553738 -960 553850 480 4 la_oenb[120]
port 423 nsew
rlabel metal2 s 557326 -960 557438 480 4 la_oenb[121]
port 424 nsew
rlabel metal2 s 560822 -960 560934 480 4 la_oenb[122]
port 425 nsew
rlabel metal2 s 564410 -960 564522 480 4 la_oenb[123]
port 426 nsew
rlabel metal2 s 567998 -960 568110 480 4 la_oenb[124]
port 427 nsew
rlabel metal2 s 571494 -960 571606 480 4 la_oenb[125]
port 428 nsew
rlabel metal2 s 575082 -960 575194 480 4 la_oenb[126]
port 429 nsew
rlabel metal2 s 578578 -960 578690 480 4 la_oenb[127]
port 430 nsew
rlabel metal2 s 170742 -960 170854 480 4 la_oenb[12]
port 431 nsew
rlabel metal2 s 174238 -960 174350 480 4 la_oenb[13]
port 432 nsew
rlabel metal2 s 177826 -960 177938 480 4 la_oenb[14]
port 433 nsew
rlabel metal2 s 181414 -960 181526 480 4 la_oenb[15]
port 434 nsew
rlabel metal2 s 184910 -960 185022 480 4 la_oenb[16]
port 435 nsew
rlabel metal2 s 188498 -960 188610 480 4 la_oenb[17]
port 436 nsew
rlabel metal2 s 191994 -960 192106 480 4 la_oenb[18]
port 437 nsew
rlabel metal2 s 195582 -960 195694 480 4 la_oenb[19]
port 438 nsew
rlabel metal2 s 131734 -960 131846 480 4 la_oenb[1]
port 439 nsew
rlabel metal2 s 199078 -960 199190 480 4 la_oenb[20]
port 440 nsew
rlabel metal2 s 202666 -960 202778 480 4 la_oenb[21]
port 441 nsew
rlabel metal2 s 206162 -960 206274 480 4 la_oenb[22]
port 442 nsew
rlabel metal2 s 209750 -960 209862 480 4 la_oenb[23]
port 443 nsew
rlabel metal2 s 213338 -960 213450 480 4 la_oenb[24]
port 444 nsew
rlabel metal2 s 216834 -960 216946 480 4 la_oenb[25]
port 445 nsew
rlabel metal2 s 220422 -960 220534 480 4 la_oenb[26]
port 446 nsew
rlabel metal2 s 223918 -960 224030 480 4 la_oenb[27]
port 447 nsew
rlabel metal2 s 227506 -960 227618 480 4 la_oenb[28]
port 448 nsew
rlabel metal2 s 231002 -960 231114 480 4 la_oenb[29]
port 449 nsew
rlabel metal2 s 135230 -960 135342 480 4 la_oenb[2]
port 450 nsew
rlabel metal2 s 234590 -960 234702 480 4 la_oenb[30]
port 451 nsew
rlabel metal2 s 238086 -960 238198 480 4 la_oenb[31]
port 452 nsew
rlabel metal2 s 241674 -960 241786 480 4 la_oenb[32]
port 453 nsew
rlabel metal2 s 245170 -960 245282 480 4 la_oenb[33]
port 454 nsew
rlabel metal2 s 248758 -960 248870 480 4 la_oenb[34]
port 455 nsew
rlabel metal2 s 252346 -960 252458 480 4 la_oenb[35]
port 456 nsew
rlabel metal2 s 255842 -960 255954 480 4 la_oenb[36]
port 457 nsew
rlabel metal2 s 259430 -960 259542 480 4 la_oenb[37]
port 458 nsew
rlabel metal2 s 262926 -960 263038 480 4 la_oenb[38]
port 459 nsew
rlabel metal2 s 266514 -960 266626 480 4 la_oenb[39]
port 460 nsew
rlabel metal2 s 138818 -960 138930 480 4 la_oenb[3]
port 461 nsew
rlabel metal2 s 270010 -960 270122 480 4 la_oenb[40]
port 462 nsew
rlabel metal2 s 273598 -960 273710 480 4 la_oenb[41]
port 463 nsew
rlabel metal2 s 277094 -960 277206 480 4 la_oenb[42]
port 464 nsew
rlabel metal2 s 280682 -960 280794 480 4 la_oenb[43]
port 465 nsew
rlabel metal2 s 284270 -960 284382 480 4 la_oenb[44]
port 466 nsew
rlabel metal2 s 287766 -960 287878 480 4 la_oenb[45]
port 467 nsew
rlabel metal2 s 291354 -960 291466 480 4 la_oenb[46]
port 468 nsew
rlabel metal2 s 294850 -960 294962 480 4 la_oenb[47]
port 469 nsew
rlabel metal2 s 298438 -960 298550 480 4 la_oenb[48]
port 470 nsew
rlabel metal2 s 301934 -960 302046 480 4 la_oenb[49]
port 471 nsew
rlabel metal2 s 142406 -960 142518 480 4 la_oenb[4]
port 472 nsew
rlabel metal2 s 305522 -960 305634 480 4 la_oenb[50]
port 473 nsew
rlabel metal2 s 309018 -960 309130 480 4 la_oenb[51]
port 474 nsew
rlabel metal2 s 312606 -960 312718 480 4 la_oenb[52]
port 475 nsew
rlabel metal2 s 316194 -960 316306 480 4 la_oenb[53]
port 476 nsew
rlabel metal2 s 319690 -960 319802 480 4 la_oenb[54]
port 477 nsew
rlabel metal2 s 323278 -960 323390 480 4 la_oenb[55]
port 478 nsew
rlabel metal2 s 326774 -960 326886 480 4 la_oenb[56]
port 479 nsew
rlabel metal2 s 330362 -960 330474 480 4 la_oenb[57]
port 480 nsew
rlabel metal2 s 333858 -960 333970 480 4 la_oenb[58]
port 481 nsew
rlabel metal2 s 337446 -960 337558 480 4 la_oenb[59]
port 482 nsew
rlabel metal2 s 145902 -960 146014 480 4 la_oenb[5]
port 483 nsew
rlabel metal2 s 340942 -960 341054 480 4 la_oenb[60]
port 484 nsew
rlabel metal2 s 344530 -960 344642 480 4 la_oenb[61]
port 485 nsew
rlabel metal2 s 348026 -960 348138 480 4 la_oenb[62]
port 486 nsew
rlabel metal2 s 351614 -960 351726 480 4 la_oenb[63]
port 487 nsew
rlabel metal2 s 355202 -960 355314 480 4 la_oenb[64]
port 488 nsew
rlabel metal2 s 358698 -960 358810 480 4 la_oenb[65]
port 489 nsew
rlabel metal2 s 362286 -960 362398 480 4 la_oenb[66]
port 490 nsew
rlabel metal2 s 365782 -960 365894 480 4 la_oenb[67]
port 491 nsew
rlabel metal2 s 369370 -960 369482 480 4 la_oenb[68]
port 492 nsew
rlabel metal2 s 372866 -960 372978 480 4 la_oenb[69]
port 493 nsew
rlabel metal2 s 149490 -960 149602 480 4 la_oenb[6]
port 494 nsew
rlabel metal2 s 376454 -960 376566 480 4 la_oenb[70]
port 495 nsew
rlabel metal2 s 379950 -960 380062 480 4 la_oenb[71]
port 496 nsew
rlabel metal2 s 383538 -960 383650 480 4 la_oenb[72]
port 497 nsew
rlabel metal2 s 387126 -960 387238 480 4 la_oenb[73]
port 498 nsew
rlabel metal2 s 390622 -960 390734 480 4 la_oenb[74]
port 499 nsew
rlabel metal2 s 394210 -960 394322 480 4 la_oenb[75]
port 500 nsew
rlabel metal2 s 397706 -960 397818 480 4 la_oenb[76]
port 501 nsew
rlabel metal2 s 401294 -960 401406 480 4 la_oenb[77]
port 502 nsew
rlabel metal2 s 404790 -960 404902 480 4 la_oenb[78]
port 503 nsew
rlabel metal2 s 408378 -960 408490 480 4 la_oenb[79]
port 504 nsew
rlabel metal2 s 152986 -960 153098 480 4 la_oenb[7]
port 505 nsew
rlabel metal2 s 411874 -960 411986 480 4 la_oenb[80]
port 506 nsew
rlabel metal2 s 415462 -960 415574 480 4 la_oenb[81]
port 507 nsew
rlabel metal2 s 418958 -960 419070 480 4 la_oenb[82]
port 508 nsew
rlabel metal2 s 422546 -960 422658 480 4 la_oenb[83]
port 509 nsew
rlabel metal2 s 426134 -960 426246 480 4 la_oenb[84]
port 510 nsew
rlabel metal2 s 429630 -960 429742 480 4 la_oenb[85]
port 511 nsew
rlabel metal2 s 433218 -960 433330 480 4 la_oenb[86]
port 512 nsew
rlabel metal2 s 436714 -960 436826 480 4 la_oenb[87]
port 513 nsew
rlabel metal2 s 440302 -960 440414 480 4 la_oenb[88]
port 514 nsew
rlabel metal2 s 443798 -960 443910 480 4 la_oenb[89]
port 515 nsew
rlabel metal2 s 156574 -960 156686 480 4 la_oenb[8]
port 516 nsew
rlabel metal2 s 447386 -960 447498 480 4 la_oenb[90]
port 517 nsew
rlabel metal2 s 450882 -960 450994 480 4 la_oenb[91]
port 518 nsew
rlabel metal2 s 454470 -960 454582 480 4 la_oenb[92]
port 519 nsew
rlabel metal2 s 458058 -960 458170 480 4 la_oenb[93]
port 520 nsew
rlabel metal2 s 461554 -960 461666 480 4 la_oenb[94]
port 521 nsew
rlabel metal2 s 465142 -960 465254 480 4 la_oenb[95]
port 522 nsew
rlabel metal2 s 468638 -960 468750 480 4 la_oenb[96]
port 523 nsew
rlabel metal2 s 472226 -960 472338 480 4 la_oenb[97]
port 524 nsew
rlabel metal2 s 475722 -960 475834 480 4 la_oenb[98]
port 525 nsew
rlabel metal2 s 479310 -960 479422 480 4 la_oenb[99]
port 526 nsew
rlabel metal2 s 160070 -960 160182 480 4 la_oenb[9]
port 527 nsew
rlabel metal2 s 579774 -960 579886 480 4 user_clock2
port 528 nsew
rlabel metal2 s 580970 -960 581082 480 4 user_irq[0]
port 529 nsew
rlabel metal2 s 582166 -960 582278 480 4 user_irq[1]
port 530 nsew
rlabel metal2 s 583362 -960 583474 480 4 user_irq[2]
port 531 nsew
rlabel metal5 s -2006 -934 585930 -314 4 vccd1
port 532 nsew
rlabel metal5 s -2966 2866 586890 3486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 38866 586890 39486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 74866 586890 75486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 110866 586890 111486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 146866 586890 147486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 182866 586890 183486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 218866 586890 219486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 254866 586890 255486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 290866 586890 291486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 326866 586890 327486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 362866 586890 363486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 398866 586890 399486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 434866 586890 435486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 470866 586890 471486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 506866 586890 507486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 542866 586890 543486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 578866 586890 579486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 614866 586890 615486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 650866 586890 651486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 686866 586890 687486 4 vccd1
port 532 nsew
rlabel metal5 s -2006 704250 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 253794 -1894 254414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 289794 -1894 290414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 325794 -1894 326414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 361794 -1894 362414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 397794 -1894 398414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 433794 -1894 434414 336000 4 vccd1
port 532 nsew
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew
rlabel metal4 s 585310 -934 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 1794 -1894 2414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 37794 -1894 38414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 73794 -1894 74414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 109794 -1894 110414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 145794 -1894 146414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 181794 -1894 182414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 217794 -1894 218414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 253794 500000 254414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 289794 500000 290414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 325794 500000 326414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 361794 500000 362414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 397794 500000 398414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 433794 500000 434414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 469794 -1894 470414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 505794 -1894 506414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 541794 -1894 542414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 577794 -1894 578414 705830 4 vccd1
port 532 nsew
rlabel metal5 s -3926 -2854 587850 -2234 4 vccd2
port 533 nsew
rlabel metal5 s -4886 6586 588810 7206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 42586 588810 43206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 78586 588810 79206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 114586 588810 115206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 150586 588810 151206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 186586 588810 187206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 222586 588810 223206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 258586 588810 259206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 294586 588810 295206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 330586 588810 331206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 366586 588810 367206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 402586 588810 403206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 438586 588810 439206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 474586 588810 475206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 510586 588810 511206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 546586 588810 547206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 582586 588810 583206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 618586 588810 619206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 654586 588810 655206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 690586 588810 691206 4 vccd2
port 533 nsew
rlabel metal5 s -3926 706170 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 257514 -3814 258134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 293514 -3814 294134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 329514 -3814 330134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 365514 -3814 366134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 401514 -3814 402134 336000 4 vccd2
port 533 nsew
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew
rlabel metal4 s 587230 -2854 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 5514 -3814 6134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 41514 -3814 42134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 77514 -3814 78134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 113514 -3814 114134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 149514 -3814 150134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 185514 -3814 186134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 221514 -3814 222134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 257514 500000 258134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 293514 500000 294134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 329514 500000 330134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 365514 500000 366134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 401514 500000 402134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 437514 -3814 438134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 473514 -3814 474134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 509514 -3814 510134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 545514 -3814 546134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 581514 -3814 582134 707750 4 vccd2
port 533 nsew
rlabel metal5 s -5846 -4774 589770 -4154 4 vdda1
port 534 nsew
rlabel metal5 s -6806 10306 590730 10926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 46306 590730 46926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 82306 590730 82926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 118306 590730 118926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 154306 590730 154926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 190306 590730 190926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 226306 590730 226926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 262306 590730 262926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 298306 590730 298926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 334306 590730 334926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 370306 590730 370926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 406306 590730 406926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 442306 590730 442926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 478306 590730 478926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 514306 590730 514926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 550306 590730 550926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 586306 590730 586926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 622306 590730 622926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 658306 590730 658926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 694306 590730 694926 4 vdda1
port 534 nsew
rlabel metal5 s -5846 708090 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 261234 -5734 261854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 297234 -5734 297854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 333234 -5734 333854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 369234 -5734 369854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 405234 -5734 405854 336000 4 vdda1
port 534 nsew
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew
rlabel metal4 s 589150 -4774 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 9234 -5734 9854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 45234 -5734 45854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 81234 -5734 81854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 117234 -5734 117854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 153234 -5734 153854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 189234 -5734 189854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 225234 -5734 225854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 261234 500000 261854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 297234 500000 297854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 333234 500000 333854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 369234 500000 369854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 405234 500000 405854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 441234 -5734 441854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 477234 -5734 477854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 513234 -5734 513854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 549234 -5734 549854 709670 4 vdda1
port 534 nsew
rlabel metal5 s -7766 -6694 591690 -6074 4 vdda2
port 535 nsew
rlabel metal5 s -8726 14026 592650 14646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 50026 592650 50646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 86026 592650 86646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 122026 592650 122646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 158026 592650 158646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 194026 592650 194646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 230026 592650 230646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 266026 592650 266646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 302026 592650 302646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 338026 592650 338646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 374026 592650 374646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 410026 592650 410646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 446026 592650 446646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 482026 592650 482646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 518026 592650 518646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 554026 592650 554646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 590026 592650 590646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 626026 592650 626646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 662026 592650 662646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 698026 592650 698646 4 vdda2
port 535 nsew
rlabel metal5 s -7766 710010 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 264954 -7654 265574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 300954 -7654 301574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 336954 -7654 337574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 372954 -7654 373574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 408954 -7654 409574 336000 4 vdda2
port 535 nsew
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew
rlabel metal4 s 591070 -6694 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 12954 -7654 13574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 48954 -7654 49574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 84954 -7654 85574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 120954 -7654 121574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 156954 -7654 157574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 192954 -7654 193574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 228954 -7654 229574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 264954 500000 265574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 300954 500000 301574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 336954 500000 337574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 372954 500000 373574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 408954 500000 409574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 444954 -7654 445574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 480954 -7654 481574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 516954 -7654 517574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 552954 -7654 553574 711590 4 vdda2
port 535 nsew
rlabel metal5 s -6806 -5734 590730 -5114 4 vssa1
port 536 nsew
rlabel metal5 s -6806 28306 590730 28926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 64306 590730 64926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 100306 590730 100926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 136306 590730 136926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 172306 590730 172926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 208306 590730 208926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 244306 590730 244926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 280306 590730 280926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 316306 590730 316926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 352306 590730 352926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 388306 590730 388926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 424306 590730 424926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 460306 590730 460926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 496306 590730 496926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 532306 590730 532926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 568306 590730 568926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 604306 590730 604926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 640306 590730 640926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 676306 590730 676926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 709050 590730 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 -5734 243854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 279234 -5734 279854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 315234 -5734 315854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 351234 -5734 351854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 387234 -5734 387854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 423234 -5734 423854 336000 4 vssa1
port 536 nsew
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew
rlabel metal4 s 27234 -5734 27854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 63234 -5734 63854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 99234 -5734 99854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 135234 -5734 135854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 171234 -5734 171854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 207234 -5734 207854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 500000 243854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 279234 500000 279854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 315234 500000 315854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 351234 500000 351854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 387234 500000 387854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 423234 500000 423854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 459234 -5734 459854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 495234 -5734 495854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 531234 -5734 531854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 567234 -5734 567854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 590110 -5734 590730 709670 4 vssa1
port 536 nsew
rlabel metal5 s -8726 -7654 592650 -7034 4 vssa2
port 537 nsew
rlabel metal5 s -8726 32026 592650 32646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 68026 592650 68646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 104026 592650 104646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 140026 592650 140646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 176026 592650 176646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 212026 592650 212646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 248026 592650 248646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 284026 592650 284646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 320026 592650 320646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 356026 592650 356646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 392026 592650 392646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 428026 592650 428646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 464026 592650 464646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 500026 592650 500646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 536026 592650 536646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 572026 592650 572646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 608026 592650 608646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 644026 592650 644646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 680026 592650 680646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 710970 592650 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 -7654 247574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 282954 -7654 283574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 318954 -7654 319574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 354954 -7654 355574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 390954 -7654 391574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 426954 -7654 427574 336000 4 vssa2
port 537 nsew
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew
rlabel metal4 s 30954 -7654 31574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 66954 -7654 67574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 102954 -7654 103574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 138954 -7654 139574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 174954 -7654 175574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 210954 -7654 211574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 500000 247574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 282954 500000 283574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 318954 500000 319574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 354954 500000 355574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 390954 500000 391574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 426954 500000 427574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 462954 -7654 463574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 498954 -7654 499574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 534954 -7654 535574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 570954 -7654 571574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 592030 -7654 592650 711590 4 vssa2
port 537 nsew
rlabel metal5 s -2966 -1894 586890 -1274 4 vssd1
port 538 nsew
rlabel metal5 s -2966 20866 586890 21486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 56866 586890 57486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 92866 586890 93486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 128866 586890 129486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 164866 586890 165486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 200866 586890 201486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 236866 586890 237486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 272866 586890 273486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 308866 586890 309486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 344866 586890 345486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 380866 586890 381486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 416866 586890 417486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 452866 586890 453486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 488866 586890 489486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 524866 586890 525486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 560866 586890 561486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 596866 586890 597486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 632866 586890 633486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 668866 586890 669486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 705210 586890 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 -1894 236414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 271794 -1894 272414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 307794 -1894 308414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 343794 -1894 344414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 379794 -1894 380414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 415794 -1894 416414 336000 4 vssd1
port 538 nsew
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew
rlabel metal4 s 19794 -1894 20414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 55794 -1894 56414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 91794 -1894 92414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 127794 -1894 128414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 163794 -1894 164414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 199794 -1894 200414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 500000 236414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 271794 500000 272414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 307794 500000 308414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 343794 500000 344414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 379794 500000 380414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 415794 500000 416414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 451794 -1894 452414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 487794 -1894 488414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 523794 -1894 524414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 559794 -1894 560414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 586270 -1894 586890 705830 4 vssd1
port 538 nsew
rlabel metal5 s -4886 -3814 588810 -3194 4 vssd2
port 539 nsew
rlabel metal5 s -4886 24586 588810 25206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 60586 588810 61206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 96586 588810 97206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 132586 588810 133206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 168586 588810 169206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 204586 588810 205206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 240586 588810 241206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 276586 588810 277206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 312586 588810 313206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 348586 588810 349206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 384586 588810 385206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 420586 588810 421206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 456586 588810 457206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 492586 588810 493206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 528586 588810 529206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 564586 588810 565206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 600586 588810 601206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 636586 588810 637206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 672586 588810 673206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 707130 588810 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 -3814 240134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 275514 -3814 276134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 311514 -3814 312134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 347514 -3814 348134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 383514 -3814 384134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 419514 -3814 420134 336000 4 vssd2
port 539 nsew
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew
rlabel metal4 s 23514 -3814 24134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 59514 -3814 60134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 95514 -3814 96134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 131514 -3814 132134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 167514 -3814 168134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 203514 -3814 204134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 500000 240134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 275514 500000 276134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 311514 500000 312134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 347514 500000 348134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 383514 500000 384134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 419514 500000 420134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 455514 -3814 456134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 491514 -3814 492134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 527514 -3814 528134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 563514 -3814 564134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 588190 -3814 588810 707750 4 vssd2
port 539 nsew
rlabel metal2 s 542 -960 654 480 4 wb_clk_i
port 540 nsew
rlabel metal2 s 1646 -960 1758 480 4 wb_rst_i
port 541 nsew
rlabel metal2 s 2842 -960 2954 480 4 wbs_ack_o
port 542 nsew
rlabel metal2 s 7626 -960 7738 480 4 wbs_adr_i[0]
port 543 nsew
rlabel metal2 s 47830 -960 47942 480 4 wbs_adr_i[10]
port 544 nsew
rlabel metal2 s 51326 -960 51438 480 4 wbs_adr_i[11]
port 545 nsew
rlabel metal2 s 54914 -960 55026 480 4 wbs_adr_i[12]
port 546 nsew
rlabel metal2 s 58410 -960 58522 480 4 wbs_adr_i[13]
port 547 nsew
rlabel metal2 s 61998 -960 62110 480 4 wbs_adr_i[14]
port 548 nsew
rlabel metal2 s 65494 -960 65606 480 4 wbs_adr_i[15]
port 549 nsew
rlabel metal2 s 69082 -960 69194 480 4 wbs_adr_i[16]
port 550 nsew
rlabel metal2 s 72578 -960 72690 480 4 wbs_adr_i[17]
port 551 nsew
rlabel metal2 s 76166 -960 76278 480 4 wbs_adr_i[18]
port 552 nsew
rlabel metal2 s 79662 -960 79774 480 4 wbs_adr_i[19]
port 553 nsew
rlabel metal2 s 12318 -960 12430 480 4 wbs_adr_i[1]
port 554 nsew
rlabel metal2 s 83250 -960 83362 480 4 wbs_adr_i[20]
port 555 nsew
rlabel metal2 s 86838 -960 86950 480 4 wbs_adr_i[21]
port 556 nsew
rlabel metal2 s 90334 -960 90446 480 4 wbs_adr_i[22]
port 557 nsew
rlabel metal2 s 93922 -960 94034 480 4 wbs_adr_i[23]
port 558 nsew
rlabel metal2 s 97418 -960 97530 480 4 wbs_adr_i[24]
port 559 nsew
rlabel metal2 s 101006 -960 101118 480 4 wbs_adr_i[25]
port 560 nsew
rlabel metal2 s 104502 -960 104614 480 4 wbs_adr_i[26]
port 561 nsew
rlabel metal2 s 108090 -960 108202 480 4 wbs_adr_i[27]
port 562 nsew
rlabel metal2 s 111586 -960 111698 480 4 wbs_adr_i[28]
port 563 nsew
rlabel metal2 s 115174 -960 115286 480 4 wbs_adr_i[29]
port 564 nsew
rlabel metal2 s 17010 -960 17122 480 4 wbs_adr_i[2]
port 565 nsew
rlabel metal2 s 118762 -960 118874 480 4 wbs_adr_i[30]
port 566 nsew
rlabel metal2 s 122258 -960 122370 480 4 wbs_adr_i[31]
port 567 nsew
rlabel metal2 s 21794 -960 21906 480 4 wbs_adr_i[3]
port 568 nsew
rlabel metal2 s 26486 -960 26598 480 4 wbs_adr_i[4]
port 569 nsew
rlabel metal2 s 30074 -960 30186 480 4 wbs_adr_i[5]
port 570 nsew
rlabel metal2 s 33570 -960 33682 480 4 wbs_adr_i[6]
port 571 nsew
rlabel metal2 s 37158 -960 37270 480 4 wbs_adr_i[7]
port 572 nsew
rlabel metal2 s 40654 -960 40766 480 4 wbs_adr_i[8]
port 573 nsew
rlabel metal2 s 44242 -960 44354 480 4 wbs_adr_i[9]
port 574 nsew
rlabel metal2 s 4038 -960 4150 480 4 wbs_cyc_i
port 575 nsew
rlabel metal2 s 8730 -960 8842 480 4 wbs_dat_i[0]
port 576 nsew
rlabel metal2 s 48934 -960 49046 480 4 wbs_dat_i[10]
port 577 nsew
rlabel metal2 s 52522 -960 52634 480 4 wbs_dat_i[11]
port 578 nsew
rlabel metal2 s 56018 -960 56130 480 4 wbs_dat_i[12]
port 579 nsew
rlabel metal2 s 59606 -960 59718 480 4 wbs_dat_i[13]
port 580 nsew
rlabel metal2 s 63194 -960 63306 480 4 wbs_dat_i[14]
port 581 nsew
rlabel metal2 s 66690 -960 66802 480 4 wbs_dat_i[15]
port 582 nsew
rlabel metal2 s 70278 -960 70390 480 4 wbs_dat_i[16]
port 583 nsew
rlabel metal2 s 73774 -960 73886 480 4 wbs_dat_i[17]
port 584 nsew
rlabel metal2 s 77362 -960 77474 480 4 wbs_dat_i[18]
port 585 nsew
rlabel metal2 s 80858 -960 80970 480 4 wbs_dat_i[19]
port 586 nsew
rlabel metal2 s 13514 -960 13626 480 4 wbs_dat_i[1]
port 587 nsew
rlabel metal2 s 84446 -960 84558 480 4 wbs_dat_i[20]
port 588 nsew
rlabel metal2 s 87942 -960 88054 480 4 wbs_dat_i[21]
port 589 nsew
rlabel metal2 s 91530 -960 91642 480 4 wbs_dat_i[22]
port 590 nsew
rlabel metal2 s 95118 -960 95230 480 4 wbs_dat_i[23]
port 591 nsew
rlabel metal2 s 98614 -960 98726 480 4 wbs_dat_i[24]
port 592 nsew
rlabel metal2 s 102202 -960 102314 480 4 wbs_dat_i[25]
port 593 nsew
rlabel metal2 s 105698 -960 105810 480 4 wbs_dat_i[26]
port 594 nsew
rlabel metal2 s 109286 -960 109398 480 4 wbs_dat_i[27]
port 595 nsew
rlabel metal2 s 112782 -960 112894 480 4 wbs_dat_i[28]
port 596 nsew
rlabel metal2 s 116370 -960 116482 480 4 wbs_dat_i[29]
port 597 nsew
rlabel metal2 s 18206 -960 18318 480 4 wbs_dat_i[2]
port 598 nsew
rlabel metal2 s 119866 -960 119978 480 4 wbs_dat_i[30]
port 599 nsew
rlabel metal2 s 123454 -960 123566 480 4 wbs_dat_i[31]
port 600 nsew
rlabel metal2 s 22990 -960 23102 480 4 wbs_dat_i[3]
port 601 nsew
rlabel metal2 s 27682 -960 27794 480 4 wbs_dat_i[4]
port 602 nsew
rlabel metal2 s 31270 -960 31382 480 4 wbs_dat_i[5]
port 603 nsew
rlabel metal2 s 34766 -960 34878 480 4 wbs_dat_i[6]
port 604 nsew
rlabel metal2 s 38354 -960 38466 480 4 wbs_dat_i[7]
port 605 nsew
rlabel metal2 s 41850 -960 41962 480 4 wbs_dat_i[8]
port 606 nsew
rlabel metal2 s 45438 -960 45550 480 4 wbs_dat_i[9]
port 607 nsew
rlabel metal2 s 9926 -960 10038 480 4 wbs_dat_o[0]
port 608 nsew
rlabel metal2 s 50130 -960 50242 480 4 wbs_dat_o[10]
port 609 nsew
rlabel metal2 s 53718 -960 53830 480 4 wbs_dat_o[11]
port 610 nsew
rlabel metal2 s 57214 -960 57326 480 4 wbs_dat_o[12]
port 611 nsew
rlabel metal2 s 60802 -960 60914 480 4 wbs_dat_o[13]
port 612 nsew
rlabel metal2 s 64298 -960 64410 480 4 wbs_dat_o[14]
port 613 nsew
rlabel metal2 s 67886 -960 67998 480 4 wbs_dat_o[15]
port 614 nsew
rlabel metal2 s 71474 -960 71586 480 4 wbs_dat_o[16]
port 615 nsew
rlabel metal2 s 74970 -960 75082 480 4 wbs_dat_o[17]
port 616 nsew
rlabel metal2 s 78558 -960 78670 480 4 wbs_dat_o[18]
port 617 nsew
rlabel metal2 s 82054 -960 82166 480 4 wbs_dat_o[19]
port 618 nsew
rlabel metal2 s 14710 -960 14822 480 4 wbs_dat_o[1]
port 619 nsew
rlabel metal2 s 85642 -960 85754 480 4 wbs_dat_o[20]
port 620 nsew
rlabel metal2 s 89138 -960 89250 480 4 wbs_dat_o[21]
port 621 nsew
rlabel metal2 s 92726 -960 92838 480 4 wbs_dat_o[22]
port 622 nsew
rlabel metal2 s 96222 -960 96334 480 4 wbs_dat_o[23]
port 623 nsew
rlabel metal2 s 99810 -960 99922 480 4 wbs_dat_o[24]
port 624 nsew
rlabel metal2 s 103306 -960 103418 480 4 wbs_dat_o[25]
port 625 nsew
rlabel metal2 s 106894 -960 107006 480 4 wbs_dat_o[26]
port 626 nsew
rlabel metal2 s 110482 -960 110594 480 4 wbs_dat_o[27]
port 627 nsew
rlabel metal2 s 113978 -960 114090 480 4 wbs_dat_o[28]
port 628 nsew
rlabel metal2 s 117566 -960 117678 480 4 wbs_dat_o[29]
port 629 nsew
rlabel metal2 s 19402 -960 19514 480 4 wbs_dat_o[2]
port 630 nsew
rlabel metal2 s 121062 -960 121174 480 4 wbs_dat_o[30]
port 631 nsew
rlabel metal2 s 124650 -960 124762 480 4 wbs_dat_o[31]
port 632 nsew
rlabel metal2 s 24186 -960 24298 480 4 wbs_dat_o[3]
port 633 nsew
rlabel metal2 s 28878 -960 28990 480 4 wbs_dat_o[4]
port 634 nsew
rlabel metal2 s 32374 -960 32486 480 4 wbs_dat_o[5]
port 635 nsew
rlabel metal2 s 35962 -960 36074 480 4 wbs_dat_o[6]
port 636 nsew
rlabel metal2 s 39550 -960 39662 480 4 wbs_dat_o[7]
port 637 nsew
rlabel metal2 s 43046 -960 43158 480 4 wbs_dat_o[8]
port 638 nsew
rlabel metal2 s 46634 -960 46746 480 4 wbs_dat_o[9]
port 639 nsew
rlabel metal2 s 11122 -960 11234 480 4 wbs_sel_i[0]
port 640 nsew
rlabel metal2 s 15906 -960 16018 480 4 wbs_sel_i[1]
port 641 nsew
rlabel metal2 s 20598 -960 20710 480 4 wbs_sel_i[2]
port 642 nsew
rlabel metal2 s 25290 -960 25402 480 4 wbs_sel_i[3]
port 643 nsew
rlabel metal2 s 5234 -960 5346 480 4 wbs_stb_i
port 644 nsew
rlabel metal2 s 6430 -960 6542 480 4 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
